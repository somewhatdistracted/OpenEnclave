../results/top.lef