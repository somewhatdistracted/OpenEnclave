`define PLAINTEXT_MODULUS 32
`define PLAINTEXT_WIDTH 5
`define DIMENSION 128
`define CIPHERTEXT_MODULUS 16777216
`define CIPHERTEXT_WIDTH 24
`define BIG_N 6425

module homomorphic_multiply_tb;

    reg clk;
    reg rst_n;
    reg [`CIPHERTEXT_WIDTH-1:0] ciphertext_entry;
    reg [`DIMENSION:0] row;
    reg ciphertext_select;
    reg en;
    wire [`CIPHERTEXT_WIDTH-1:0] result;
    reg [`CIPHERTEXT_WIDTH-1:0] expected;

    always #10 clk = ~clk;

    homomorphic_multiply #(
        .PLAINTEXT_MODULUS(`PLAINTEXT_MODULUS),
        .PLAINTEXT_WIDTH(`PLAINTEXT_WIDTH),
        .CIPHERTEXT_MODULUS(`CIPHERTEXT_MODULUS),
        .CIPHERTEXT_WIDTH(`CIPHERTEXT_WIDTH),
        .DIMENSION(`DIMENSION),
        .BIG_N(`BIG_N)
    ) homomorphic_inst (
        .clk(clk),
        .rst_n(rst_n),
        .ciphertext_entry(ciphertext_entry),
        .row(row),
        .ciphertext_select(ciphertext_select),
        .en(en),
        .result_partial(result)
    );

    initial begin
        clk = 0;
        ciphertext_select = 0;
        row = 0;
        ciphertext_entry = 0;

en=0;
rst_n=0;
#100;
rst_n=1;
#100;
en=1;
ciphertext_select = 0;
row = 0;
ciphertext_entry =8556363;
#20;
row = 1;
ciphertext_entry =11084185;
#20;
row = 2;
ciphertext_entry =10350093;
#20;
row = 3;
ciphertext_entry =8355122;
#20;
row = 4;
ciphertext_entry =763708;
#20;
row = 5;
ciphertext_entry =15427112;
#20;
row = 6;
ciphertext_entry =10902113;
#20;
row = 7;
ciphertext_entry =9960714;
#20;
row = 8;
ciphertext_entry =3119218;
#20;
row = 9;
ciphertext_entry =9531090;
#20;
row = 10;
ciphertext_entry =9386273;
#20;
row = 11;
ciphertext_entry =1133811;
#20;
row = 12;
ciphertext_entry =15639104;
#20;
row = 13;
ciphertext_entry =10781349;
#20;
row = 14;
ciphertext_entry =3034581;
#20;
row = 15;
ciphertext_entry =12675627;
#20;
row = 16;
ciphertext_entry =862728;
#20;
row = 17;
ciphertext_entry =13626759;
#20;
row = 18;
ciphertext_entry =6931480;
#20;
row = 19;
ciphertext_entry =5507229;
#20;
row = 20;
ciphertext_entry =1765353;
#20;
row = 21;
ciphertext_entry =5562099;
#20;
row = 22;
ciphertext_entry =668709;
#20;
row = 23;
ciphertext_entry =9330992;
#20;
row = 24;
ciphertext_entry =16159103;
#20;
row = 25;
ciphertext_entry =11150655;
#20;
row = 26;
ciphertext_entry =13827912;
#20;
row = 27;
ciphertext_entry =5933645;
#20;
row = 28;
ciphertext_entry =5503615;
#20;
row = 29;
ciphertext_entry =4114011;
#20;
row = 30;
ciphertext_entry =4279505;
#20;
row = 31;
ciphertext_entry =8545352;
#20;
row = 32;
ciphertext_entry =823104;
#20;
row = 33;
ciphertext_entry =8297742;
#20;
row = 34;
ciphertext_entry =7419884;
#20;
row = 35;
ciphertext_entry =15194888;
#20;
row = 36;
ciphertext_entry =15658189;
#20;
row = 37;
ciphertext_entry =11920927;
#20;
row = 38;
ciphertext_entry =4689677;
#20;
row = 39;
ciphertext_entry =8034167;
#20;
row = 40;
ciphertext_entry =14666369;
#20;
row = 41;
ciphertext_entry =8166148;
#20;
row = 42;
ciphertext_entry =9737606;
#20;
row = 43;
ciphertext_entry =10954692;
#20;
row = 44;
ciphertext_entry =7480455;
#20;
row = 45;
ciphertext_entry =8874230;
#20;
row = 46;
ciphertext_entry =6095977;
#20;
row = 47;
ciphertext_entry =4117651;
#20;
row = 48;
ciphertext_entry =6777835;
#20;
row = 49;
ciphertext_entry =16680523;
#20;
row = 50;
ciphertext_entry =12766457;
#20;
row = 51;
ciphertext_entry =13675935;
#20;
row = 52;
ciphertext_entry =3960481;
#20;
row = 53;
ciphertext_entry =9969573;
#20;
row = 54;
ciphertext_entry =14919880;
#20;
row = 55;
ciphertext_entry =12288347;
#20;
row = 56;
ciphertext_entry =3414621;
#20;
row = 57;
ciphertext_entry =9023805;
#20;
row = 58;
ciphertext_entry =3410032;
#20;
row = 59;
ciphertext_entry =11074170;
#20;
row = 60;
ciphertext_entry =376918;
#20;
row = 61;
ciphertext_entry =11542885;
#20;
row = 62;
ciphertext_entry =1023003;
#20;
row = 63;
ciphertext_entry =9043181;
#20;
row = 64;
ciphertext_entry =7691292;
#20;
row = 65;
ciphertext_entry =6461981;
#20;
row = 66;
ciphertext_entry =8795965;
#20;
row = 67;
ciphertext_entry =10341406;
#20;
row = 68;
ciphertext_entry =16517278;
#20;
row = 69;
ciphertext_entry =1722607;
#20;
row = 70;
ciphertext_entry =13080491;
#20;
row = 71;
ciphertext_entry =13714605;
#20;
row = 72;
ciphertext_entry =4780423;
#20;
row = 73;
ciphertext_entry =1341041;
#20;
row = 74;
ciphertext_entry =40318;
#20;
row = 75;
ciphertext_entry =8839059;
#20;
row = 76;
ciphertext_entry =11605193;
#20;
row = 77;
ciphertext_entry =7682761;
#20;
row = 78;
ciphertext_entry =14244716;
#20;
row = 79;
ciphertext_entry =3211433;
#20;
row = 80;
ciphertext_entry =16047061;
#20;
row = 81;
ciphertext_entry =16641399;
#20;
row = 82;
ciphertext_entry =12820358;
#20;
row = 83;
ciphertext_entry =14579095;
#20;
row = 84;
ciphertext_entry =12861938;
#20;
row = 85;
ciphertext_entry =9826068;
#20;
row = 86;
ciphertext_entry =4720495;
#20;
row = 87;
ciphertext_entry =1440193;
#20;
row = 88;
ciphertext_entry =7327947;
#20;
row = 89;
ciphertext_entry =14674863;
#20;
row = 90;
ciphertext_entry =1119017;
#20;
row = 91;
ciphertext_entry =5465961;
#20;
row = 92;
ciphertext_entry =6478166;
#20;
row = 93;
ciphertext_entry =9361734;
#20;
row = 94;
ciphertext_entry =3400125;
#20;
row = 95;
ciphertext_entry =8991956;
#20;
row = 96;
ciphertext_entry =13846085;
#20;
row = 97;
ciphertext_entry =8343959;
#20;
row = 98;
ciphertext_entry =10039498;
#20;
row = 99;
ciphertext_entry =11959258;
#20;
row = 100;
ciphertext_entry =2623572;
#20;
row = 101;
ciphertext_entry =1809431;
#20;
row = 102;
ciphertext_entry =11886750;
#20;
row = 103;
ciphertext_entry =8466456;
#20;
row = 104;
ciphertext_entry =3612884;
#20;
row = 105;
ciphertext_entry =5634223;
#20;
row = 106;
ciphertext_entry =5049772;
#20;
row = 107;
ciphertext_entry =15597315;
#20;
row = 108;
ciphertext_entry =1313191;
#20;
row = 109;
ciphertext_entry =6705617;
#20;
row = 110;
ciphertext_entry =14354095;
#20;
row = 111;
ciphertext_entry =495375;
#20;
row = 112;
ciphertext_entry =5246060;
#20;
row = 113;
ciphertext_entry =14913974;
#20;
row = 114;
ciphertext_entry =1314112;
#20;
row = 115;
ciphertext_entry =13016199;
#20;
row = 116;
ciphertext_entry =16253714;
#20;
row = 117;
ciphertext_entry =1358191;
#20;
row = 118;
ciphertext_entry =3129399;
#20;
row = 119;
ciphertext_entry =10736031;
#20;
row = 120;
ciphertext_entry =11453872;
#20;
row = 121;
ciphertext_entry =13447415;
#20;
row = 122;
ciphertext_entry =15741607;
#20;
row = 123;
ciphertext_entry =2605416;
#20;
row = 124;
ciphertext_entry =6406665;
#20;
row = 125;
ciphertext_entry =10738357;
#20;
row = 126;
ciphertext_entry =11461538;
#20;
row = 127;
ciphertext_entry =7666522;
#20;
row = 128;
ciphertext_entry =6339490;
#20;
ciphertext_select = 1;
row = 0;
ciphertext_entry =8556363;
#20;
$display("Result = %d", result); assert(result ==8544600);
row = 1;
ciphertext_entry =11084185;
#20;
$display("Result = %d", result); assert(result ==2066817);
row = 2;
ciphertext_entry =10350093;
#20;
$display("Result = %d", result); assert(result ==8417256);
row = 3;
ciphertext_entry =8355122;
#20;
$display("Result = %d", result); assert(result ==16360709);
row = 4;
ciphertext_entry =763708;
#20;
$display("Result = %d", result); assert(result ==1308439);
row = 5;
ciphertext_entry =15427112;
#20;
$display("Result = %d", result); assert(result ==12483703);
row = 6;
ciphertext_entry =10902113;
#20;
$display("Result = %d", result); assert(result ==12798281);
row = 7;
ciphertext_entry =9960714;
#20;
$display("Result = %d", result); assert(result ==12082981);
row = 8;
ciphertext_entry =3119218;
#20;
$display("Result = %d", result); assert(result ==9109583);
row = 9;
ciphertext_entry =9531090;
#20;
$display("Result = %d", result); assert(result ==1184048);
row = 10;
ciphertext_entry =9386273;
#20;
$display("Result = %d", result); assert(result ==13992875);
row = 11;
ciphertext_entry =1133811;
#20;
$display("Result = %d", result); assert(result ==8539957);
row = 12;
ciphertext_entry =15639104;
#20;
$display("Result = %d", result); assert(result ==3415234);
row = 13;
ciphertext_entry =10781349;
#20;
$display("Result = %d", result); assert(result ==4707799);
row = 14;
ciphertext_entry =3034581;
#20;
$display("Result = %d", result); assert(result ==16717603);
row = 15;
ciphertext_entry =12675627;
#20;
$display("Result = %d", result); assert(result ==8374105);
row = 16;
ciphertext_entry =862728;
#20;
$display("Result = %d", result); assert(result ==13211720);
row = 17;
ciphertext_entry =13626759;
#20;
$display("Result = %d", result); assert(result ==12749984);
row = 18;
ciphertext_entry =6931480;
#20;
$display("Result = %d", result); assert(result ==5120547);
row = 19;
ciphertext_entry =5507229;
#20;
$display("Result = %d", result); assert(result ==15365386);
row = 20;
ciphertext_entry =1765353;
#20;
$display("Result = %d", result); assert(result ==12064182);
row = 21;
ciphertext_entry =5562099;
#20;
$display("Result = %d", result); assert(result ==4488388);
row = 22;
ciphertext_entry =668709;
#20;
$display("Result = %d", result); assert(result ==12002151);
row = 23;
ciphertext_entry =9330992;
#20;
$display("Result = %d", result); assert(result ==8312025);
row = 24;
ciphertext_entry =16159103;
#20;
$display("Result = %d", result); assert(result ==14551565);
row = 25;
ciphertext_entry =11150655;
#20;
$display("Result = %d", result); assert(result ==13449651);
row = 26;
ciphertext_entry =13827912;
#20;
$display("Result = %d", result); assert(result ==5658855);
row = 27;
ciphertext_entry =5933645;
#20;
$display("Result = %d", result); assert(result ==1647430);
row = 28;
ciphertext_entry =5503615;
#20;
$display("Result = %d", result); assert(result ==3575174);
row = 29;
ciphertext_entry =4114011;
#20;
$display("Result = %d", result); assert(result ==4379309);
row = 30;
ciphertext_entry =4279505;
#20;
$display("Result = %d", result); assert(result ==10680073);
row = 31;
ciphertext_entry =8545352;
#20;
$display("Result = %d", result); assert(result ==1558222);
row = 32;
ciphertext_entry =823104;
#20;
$display("Result = %d", result); assert(result ==4127660);
row = 33;
ciphertext_entry =8297742;
#20;
$display("Result = %d", result); assert(result ==2433889);
row = 34;
ciphertext_entry =7419884;
#20;
$display("Result = %d", result); assert(result ==7772752);
row = 35;
ciphertext_entry =15194888;
#20;
$display("Result = %d", result); assert(result ==3165750);
row = 36;
ciphertext_entry =15658189;
#20;
$display("Result = %d", result); assert(result ==6781756);
row = 37;
ciphertext_entry =11920927;
#20;
$display("Result = %d", result); assert(result ==12905795);
row = 38;
ciphertext_entry =4689677;
#20;
$display("Result = %d", result); assert(result ==8991667);
row = 39;
ciphertext_entry =8034167;
#20;
$display("Result = %d", result); assert(result ==12680115);
row = 40;
ciphertext_entry =14666369;
#20;
$display("Result = %d", result); assert(result ==15016204);
row = 41;
ciphertext_entry =8166148;
#20;
$display("Result = %d", result); assert(result ==5675977);
row = 42;
ciphertext_entry =9737606;
#20;
$display("Result = %d", result); assert(result ==14778561);
row = 43;
ciphertext_entry =10954692;
#20;
$display("Result = %d", result); assert(result ==3372161);
row = 44;
ciphertext_entry =7480455;
#20;
$display("Result = %d", result); assert(result ==13726329);
row = 45;
ciphertext_entry =8874230;
#20;
$display("Result = %d", result); assert(result ==10039854);
row = 46;
ciphertext_entry =6095977;
#20;
$display("Result = %d", result); assert(result ==3759430);
row = 47;
ciphertext_entry =4117651;
#20;
$display("Result = %d", result); assert(result ==4118295);
row = 48;
ciphertext_entry =6777835;
#20;
$display("Result = %d", result); assert(result ==13273504);
row = 49;
ciphertext_entry =16680523;
#20;
$display("Result = %d", result); assert(result ==5412875);
row = 50;
ciphertext_entry =12766457;
#20;
$display("Result = %d", result); assert(result ==5894253);
row = 51;
ciphertext_entry =13675935;
#20;
$display("Result = %d", result); assert(result ==4259791);
row = 52;
ciphertext_entry =3960481;
#20;
$display("Result = %d", result); assert(result ==9257756);
row = 53;
ciphertext_entry =9969573;
#20;
$display("Result = %d", result); assert(result ==7071757);
row = 54;
ciphertext_entry =14919880;
#20;
$display("Result = %d", result); assert(result ==8668287);
row = 55;
ciphertext_entry =12288347;
#20;
$display("Result = %d", result); assert(result ==11636956);
row = 56;
ciphertext_entry =3414621;
#20;
$display("Result = %d", result); assert(result ==4765474);
row = 57;
ciphertext_entry =9023805;
#20;
$display("Result = %d", result); assert(result ==14173266);
row = 58;
ciphertext_entry =3410032;
#20;
$display("Result = %d", result); assert(result ==765883);
row = 59;
ciphertext_entry =11074170;
#20;
$display("Result = %d", result); assert(result ==661820);
row = 60;
ciphertext_entry =376918;
#20;
$display("Result = %d", result); assert(result ==10522777);
row = 61;
ciphertext_entry =11542885;
#20;
$display("Result = %d", result); assert(result ==15683015);
row = 62;
ciphertext_entry =1023003;
#20;
$display("Result = %d", result); assert(result ==3507609);
row = 63;
ciphertext_entry =9043181;
#20;
$display("Result = %d", result); assert(result ==3014743);
row = 64;
ciphertext_entry =7691292;
#20;
$display("Result = %d", result); assert(result ==3233504);
row = 65;
ciphertext_entry =6461981;
#20;
$display("Result = %d", result); assert(result ==8360821);
row = 66;
ciphertext_entry =8795965;
#20;
$display("Result = %d", result); assert(result ==4633209);
row = 67;
ciphertext_entry =10341406;
#20;
$display("Result = %d", result); assert(result ==7330303);
row = 68;
ciphertext_entry =16517278;
#20;
$display("Result = %d", result); assert(result ==4147118);
row = 69;
ciphertext_entry =1722607;
#20;
$display("Result = %d", result); assert(result ==766751);
row = 70;
ciphertext_entry =13080491;
#20;
$display("Result = %d", result); assert(result ==11391851);
row = 71;
ciphertext_entry =13714605;
#20;
$display("Result = %d", result); assert(result ==14236841);
row = 72;
ciphertext_entry =4780423;
#20;
$display("Result = %d", result); assert(result ==1653487);
row = 73;
ciphertext_entry =1341041;
#20;
$display("Result = %d", result); assert(result ==12780568);
row = 74;
ciphertext_entry =40318;
#20;
$display("Result = %d", result); assert(result ==15920976);
row = 75;
ciphertext_entry =8839059;
#20;
$display("Result = %d", result); assert(result ==6127868);
row = 76;
ciphertext_entry =11605193;
#20;
$display("Result = %d", result); assert(result ==1506914);
row = 77;
ciphertext_entry =7682761;
#20;
$display("Result = %d", result); assert(result ==3839977);
row = 78;
ciphertext_entry =14244716;
#20;
$display("Result = %d", result); assert(result ==13904296);
row = 79;
ciphertext_entry =3211433;
#20;
$display("Result = %d", result); assert(result ==7874995);
row = 80;
ciphertext_entry =16047061;
#20;
$display("Result = %d", result); assert(result ==9411483);
row = 81;
ciphertext_entry =16641399;
#20;
$display("Result = %d", result); assert(result ==5706485);
row = 82;
ciphertext_entry =12820358;
#20;
$display("Result = %d", result); assert(result ==375228);
row = 83;
ciphertext_entry =14579095;
#20;
$display("Result = %d", result); assert(result ==3638548);
row = 84;
ciphertext_entry =12861938;
#20;
$display("Result = %d", result); assert(result ==12860428);
row = 85;
ciphertext_entry =9826068;
#20;
$display("Result = %d", result); assert(result ==7791853);
row = 86;
ciphertext_entry =4720495;
#20;
$display("Result = %d", result); assert(result ==9422441);
row = 87;
ciphertext_entry =1440193;
#20;
$display("Result = %d", result); assert(result ==5177371);
row = 88;
ciphertext_entry =7327947;
#20;
$display("Result = %d", result); assert(result ==15655850);
row = 89;
ciphertext_entry =14674863;
#20;
$display("Result = %d", result); assert(result ==1928673);
row = 90;
ciphertext_entry =1119017;
#20;
$display("Result = %d", result); assert(result ==6165403);
row = 91;
ciphertext_entry =5465961;
#20;
$display("Result = %d", result); assert(result ==6694274);
row = 92;
ciphertext_entry =6478166;
#20;
$display("Result = %d", result); assert(result ==2818723);
row = 93;
ciphertext_entry =9361734;
#20;
$display("Result = %d", result); assert(result ==16772694);
row = 94;
ciphertext_entry =3400125;
#20;
$display("Result = %d", result); assert(result ==10344596);
row = 95;
ciphertext_entry =8991956;
#20;
$display("Result = %d", result); assert(result ==608998);
row = 96;
ciphertext_entry =13846085;
#20;
$display("Result = %d", result); assert(result ==8882830);
row = 97;
ciphertext_entry =8343959;
#20;
$display("Result = %d", result); assert(result ==13008054);
row = 98;
ciphertext_entry =10039498;
#20;
$display("Result = %d", result); assert(result ==3087721);
row = 99;
ciphertext_entry =11959258;
#20;
$display("Result = %d", result); assert(result ==13670093);
row = 100;
ciphertext_entry =2623572;
#20;
$display("Result = %d", result); assert(result ==12628045);
row = 101;
ciphertext_entry =1809431;
#20;
$display("Result = %d", result); assert(result ==14830222);
row = 102;
ciphertext_entry =11886750;
#20;
$display("Result = %d", result); assert(result ==4201307);
row = 103;
ciphertext_entry =8466456;
#20;
$display("Result = %d", result); assert(result ==5894881);
row = 104;
ciphertext_entry =3612884;
#20;
$display("Result = %d", result); assert(result ==5810988);
row = 105;
ciphertext_entry =5634223;
#20;
$display("Result = %d", result); assert(result ==4944822);
row = 106;
ciphertext_entry =5049772;
#20;
$display("Result = %d", result); assert(result ==13390244);
row = 107;
ciphertext_entry =15597315;
#20;
$display("Result = %d", result); assert(result ==5116583);
row = 108;
ciphertext_entry =1313191;
#20;
$display("Result = %d", result); assert(result ==4758959);
row = 109;
ciphertext_entry =6705617;
#20;
$display("Result = %d", result); assert(result ==327719);
row = 110;
ciphertext_entry =14354095;
#20;
$display("Result = %d", result); assert(result ==16496739);
row = 111;
ciphertext_entry =495375;
#20;
$display("Result = %d", result); assert(result ==7501080);
row = 112;
ciphertext_entry =5246060;
#20;
$display("Result = %d", result); assert(result ==8105139);
row = 113;
ciphertext_entry =14913974;
#20;
$display("Result = %d", result); assert(result ==14996431);
row = 114;
ciphertext_entry =1314112;
#20;
$display("Result = %d", result); assert(result ==12576285);
row = 115;
ciphertext_entry =13016199;
#20;
$display("Result = %d", result); assert(result ==2377009);
row = 116;
ciphertext_entry =16253714;
#20;
$display("Result = %d", result); assert(result ==8730106);
row = 117;
ciphertext_entry =1358191;
#20;
$display("Result = %d", result); assert(result ==8850045);
row = 118;
ciphertext_entry =3129399;
#20;
$display("Result = %d", result); assert(result ==3677805);
row = 119;
ciphertext_entry =10736031;
#20;
$display("Result = %d", result); assert(result ==2817151);
row = 120;
ciphertext_entry =11453872;
#20;
$display("Result = %d", result); assert(result ==15072855);
row = 121;
ciphertext_entry =13447415;
#20;
$display("Result = %d", result); assert(result ==1070205);
row = 122;
ciphertext_entry =15741607;
#20;
$display("Result = %d", result); assert(result ==7266241);
row = 123;
ciphertext_entry =2605416;
#20;
$display("Result = %d", result); assert(result ==9793034);
row = 124;
ciphertext_entry =6406665;
#20;
$display("Result = %d", result); assert(result ==12141613);
row = 125;
ciphertext_entry =10738357;
#20;
$display("Result = %d", result); assert(result ==3905558);
row = 126;
ciphertext_entry =11461538;
#20;
$display("Result = %d", result); assert(result ==10395340);
row = 127;
ciphertext_entry =7666522;
#20;
$display("Result = %d", result); assert(result ==16707784);
row = 128;
ciphertext_entry =6339490;
#20;
$display("Result = %d", result); assert(result ==3090487);
ciphertext_select = 0;
row = 129;
#20;
$display("Result = %d", result); assert(result ==12682043);
row = 130;
#20;
$display("Result = %d", result); assert(result ==1497847);
row = 131;
#20;
$display("Result = %d", result); assert(result ==13816709);
row = 132;
#20;
$display("Result = %d", result); assert(result ==12348766);
row = 133;
#20;
$display("Result = %d", result); assert(result ==8782959);
row = 134;
#20;
$display("Result = %d", result); assert(result ==14784315);
row = 135;
#20;
$display("Result = %d", result); assert(result ==9466835);
row = 136;
#20;
$display("Result = %d", result); assert(result ==9370296);
row = 137;
#20;
$display("Result = %d", result); assert(result ==10597516);
row = 138;
#20;
$display("Result = %d", result); assert(result ==1219595);
row = 139;
#20;
$display("Result = %d", result); assert(result ==10723135);
row = 140;
#20;
$display("Result = %d", result); assert(result ==3701223);
row = 141;
#20;
$display("Result = %d", result); assert(result ==916880);
row = 142;
#20;
$display("Result = %d", result); assert(result ==2650257);
row = 143;
#20;
$display("Result = %d", result); assert(result ==2826009);
row = 144;
#20;
$display("Result = %d", result); assert(result ==10615178);
row = 145;
#20;
$display("Result = %d", result); assert(result ==5054944);
row = 146;
#20;
$display("Result = %d", result); assert(result ==11565531);
row = 147;
#20;
$display("Result = %d", result); assert(result ==11289913);
row = 148;
#20;
$display("Result = %d", result); assert(result ==13294317);
row = 149;
#20;
$display("Result = %d", result); assert(result ==15468997);
row = 150;
#20;
$display("Result = %d", result); assert(result ==16255304);
row = 151;
#20;
$display("Result = %d", result); assert(result ==5361107);
row = 152;
#20;
$display("Result = %d", result); assert(result ==1534719);
row = 153;
#20;
$display("Result = %d", result); assert(result ==5071228);
row = 154;
#20;
$display("Result = %d", result); assert(result ==4909424);
row = 155;
#20;
$display("Result = %d", result); assert(result ==7876266);
row = 156;
#20;
$display("Result = %d", result); assert(result ==12521215);
row = 157;
#20;
$display("Result = %d", result); assert(result ==2100746);
row = 158;
#20;
$display("Result = %d", result); assert(result ==6112368);
row = 159;
#20;
$display("Result = %d", result); assert(result ==7643728);
row = 160;
#20;
$display("Result = %d", result); assert(result ==13247327);
row = 161;
#20;
$display("Result = %d", result); assert(result ==6497211);
row = 162;
#20;
$display("Result = %d", result); assert(result ==10919763);
row = 163;
#20;
$display("Result = %d", result); assert(result ==12892768);
row = 164;
#20;
$display("Result = %d", result); assert(result ==7070970);
row = 165;
#20;
$display("Result = %d", result); assert(result ==15841687);
row = 166;
#20;
$display("Result = %d", result); assert(result ==10172497);
row = 167;
#20;
$display("Result = %d", result); assert(result ==6018418);
row = 168;
#20;
$display("Result = %d", result); assert(result ==6134552);
row = 169;
#20;
$display("Result = %d", result); assert(result ==10560854);
row = 170;
#20;
$display("Result = %d", result); assert(result ==12440347);
row = 171;
#20;
$display("Result = %d", result); assert(result ==6673196);
row = 172;
#20;
$display("Result = %d", result); assert(result ==6977425);
row = 173;
#20;
$display("Result = %d", result); assert(result ==14319779);
row = 174;
#20;
$display("Result = %d", result); assert(result ==13715845);
row = 175;
#20;
$display("Result = %d", result); assert(result ==3699946);
row = 176;
#20;
$display("Result = %d", result); assert(result ==15577029);
row = 177;
#20;
$display("Result = %d", result); assert(result ==14034900);
row = 178;
#20;
$display("Result = %d", result); assert(result ==2082752);
row = 179;
#20;
$display("Result = %d", result); assert(result ==15568085);
row = 180;
#20;
$display("Result = %d", result); assert(result ==4529002);
row = 181;
#20;
$display("Result = %d", result); assert(result ==11049272);
row = 182;
#20;
$display("Result = %d", result); assert(result ==5927889);
row = 183;
#20;
$display("Result = %d", result); assert(result ==3418127);
row = 184;
#20;
$display("Result = %d", result); assert(result ==415995);
row = 185;
#20;
$display("Result = %d", result); assert(result ==13621569);
row = 186;
#20;
$display("Result = %d", result); assert(result ==14894220);
row = 187;
#20;
$display("Result = %d", result); assert(result ==3396197);
row = 188;
#20;
$display("Result = %d", result); assert(result ==1856610);
row = 189;
#20;
$display("Result = %d", result); assert(result ==268594);
row = 190;
#20;
$display("Result = %d", result); assert(result ==10975518);
row = 191;
#20;
$display("Result = %d", result); assert(result ==892583);
row = 192;
#20;
$display("Result = %d", result); assert(result ==6751125);
row = 193;
#20;
$display("Result = %d", result); assert(result ==4335290);
row = 194;
#20;
$display("Result = %d", result); assert(result ==11127077);
row = 195;
#20;
$display("Result = %d", result); assert(result ==15061498);
row = 196;
#20;
$display("Result = %d", result); assert(result ==2126234);
row = 197;
#20;
$display("Result = %d", result); assert(result ==10180381);
row = 198;
#20;
$display("Result = %d", result); assert(result ==13449814);
row = 199;
#20;
$display("Result = %d", result); assert(result ==16071542);
row = 200;
#20;
$display("Result = %d", result); assert(result ==2161);
row = 201;
#20;
$display("Result = %d", result); assert(result ==8504769);
row = 202;
#20;
$display("Result = %d", result); assert(result ==16256996);
row = 203;
#20;
$display("Result = %d", result); assert(result ==3746325);
row = 204;
#20;
$display("Result = %d", result); assert(result ==1436921);
row = 205;
#20;
$display("Result = %d", result); assert(result ==16570905);
row = 206;
#20;
$display("Result = %d", result); assert(result ==424834);
row = 207;
#20;
$display("Result = %d", result); assert(result ==14373293);
row = 208;
#20;
$display("Result = %d", result); assert(result ==7688631);
row = 209;
#20;
$display("Result = %d", result); assert(result ==1339487);
row = 210;
#20;
$display("Result = %d", result); assert(result ==15872898);
row = 211;
#20;
$display("Result = %d", result); assert(result ==10712605);
row = 212;
#20;
$display("Result = %d", result); assert(result ==15007067);
row = 213;
#20;
$display("Result = %d", result); assert(result ==2023407);
row = 214;
#20;
$display("Result = %d", result); assert(result ==8503622);
row = 215;
#20;
$display("Result = %d", result); assert(result ==11023009);
row = 216;
#20;
$display("Result = %d", result); assert(result ==11557895);
row = 217;
#20;
$display("Result = %d", result); assert(result ==15856772);
row = 218;
#20;
$display("Result = %d", result); assert(result ==14994244);
row = 219;
#20;
$display("Result = %d", result); assert(result ==15655135);
row = 220;
#20;
$display("Result = %d", result); assert(result ==10349385);
row = 221;
#20;
$display("Result = %d", result); assert(result ==2733556);
row = 222;
#20;
$display("Result = %d", result); assert(result ==14921664);
row = 223;
#20;
$display("Result = %d", result); assert(result ==1631304);
row = 224;
#20;
$display("Result = %d", result); assert(result ==15972235);
row = 225;
#20;
$display("Result = %d", result); assert(result ==2515828);
row = 226;
#20;
$display("Result = %d", result); assert(result ==3305228);
row = 227;
#20;
$display("Result = %d", result); assert(result ==13304433);
row = 228;
#20;
$display("Result = %d", result); assert(result ==8737794);
row = 229;
#20;
$display("Result = %d", result); assert(result ==7007382);
row = 230;
#20;
$display("Result = %d", result); assert(result ==1289670);
row = 231;
#20;
$display("Result = %d", result); assert(result ==4832969);
row = 232;
#20;
$display("Result = %d", result); assert(result ==9126504);
row = 233;
#20;
$display("Result = %d", result); assert(result ==1641758);
row = 234;
#20;
$display("Result = %d", result); assert(result ==7181373);
row = 235;
#20;
$display("Result = %d", result); assert(result ==13662790);
row = 236;
#20;
$display("Result = %d", result); assert(result ==326917);
row = 237;
#20;
$display("Result = %d", result); assert(result ==132619);
row = 238;
#20;
$display("Result = %d", result); assert(result ==47338);
row = 239;
#20;
$display("Result = %d", result); assert(result ==8378603);
row = 240;
#20;
$display("Result = %d", result); assert(result ==10406634);
row = 241;
#20;
$display("Result = %d", result); assert(result ==12613883);
row = 242;
#20;
$display("Result = %d", result); assert(result ==11842396);
row = 243;
#20;
$display("Result = %d", result); assert(result ==10128190);
row = 244;
#20;
$display("Result = %d", result); assert(result ==2807919);
row = 245;
#20;
$display("Result = %d", result); assert(result ==13925940);
row = 246;
#20;
$display("Result = %d", result); assert(result ==3523700);
row = 247;
#20;
$display("Result = %d", result); assert(result ==11747900);
row = 248;
#20;
$display("Result = %d", result); assert(result ==13243710);
row = 249;
#20;
$display("Result = %d", result); assert(result ==16195784);
row = 250;
#20;
$display("Result = %d", result); assert(result ==7269199);
row = 251;
#20;
$display("Result = %d", result); assert(result ==3523697);
row = 252;
#20;
$display("Result = %d", result); assert(result ==6684504);
row = 253;
#20;
$display("Result = %d", result); assert(result ==13210623);
row = 254;
#20;
$display("Result = %d", result); assert(result ==12912200);
row = 255;
#20;
$display("Result = %d", result); assert(result ==12581128);
row = 256;
#20;
$display("Result = %d", result); assert(result ==13168706);

$finish;
end
endmodule