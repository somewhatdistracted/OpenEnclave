`define PLAINTEXT_MODULUS 32
`define PLAINTEXT_WIDTH 5
`define DIMENSION 128
`define CIPHERTEXT_MODULUS 16777216
`define CIPHERTEXT_WIDTH 24
`define BIG_N 6425

module encrypt_tb_full;

    reg clk;
    reg rst_n;

    reg go;
    reg [`PLAINTEXT_WIDTH-1:0] plaintext;
    reg [`CIPHERTEXT_WIDTH-1:0] publickey_row [`BIG_N-1:0];
    reg [`BIG_N-1:0] noise_select;
    reg [`DIMENSION:0] row;
    reg [`CIPHERTEXT_WIDTH-1:0] ciphertext;
    reg [`CIPHERTEXT_WIDTH-1:0] expected;

    always #10 clk = ~clk;

    encrypt #(
        .PLAINTEXT_MODULUS(`PLAINTEXT_MODULUS),
        .PLAINTEXT_WIDTH(`PLAINTEXT_WIDTH),
        .CIPHERTEXT_MODULUS(`CIPHERTEXT_MODULUS),
        .CIPHERTEXT_WIDTH(`CIPHERTEXT_WIDTH),
        .DIMENSION(`DIMENSION),
        .BIG_N(`BIG_N)
    ) encrypt_inst (
        .clk(clk),
        .rst_n(rst_n),
        .plaintext(plaintext),
        .publickey_row(publickey_row),
        .noise_select(noise_select),
        .row(row),
        .ciphertext(ciphertext)
    );

    initial begin
        row = 0;
        rst_n = 1;
        go = 0;
        plaintext = 0;
        noise_select = 0;

#20

publickey_row[0] = `CIPHERTEXT_WIDTH'd1464055;
publickey_row[1] = `CIPHERTEXT_WIDTH'd1141353;
publickey_row[2] = `CIPHERTEXT_WIDTH'd14365671;
publickey_row[3] = `CIPHERTEXT_WIDTH'd8462756;
publickey_row[4] = `CIPHERTEXT_WIDTH'd13501708;
publickey_row[5] = `CIPHERTEXT_WIDTH'd7418709;
publickey_row[6] = `CIPHERTEXT_WIDTH'd14817999;
publickey_row[7] = `CIPHERTEXT_WIDTH'd15301565;
publickey_row[8] = `CIPHERTEXT_WIDTH'd2898572;
publickey_row[9] = `CIPHERTEXT_WIDTH'd6108250;
publickey_row[10] = `CIPHERTEXT_WIDTH'd9087247;
publickey_row[11] = `CIPHERTEXT_WIDTH'd14817859;
publickey_row[12] = `CIPHERTEXT_WIDTH'd14537421;
publickey_row[13] = `CIPHERTEXT_WIDTH'd4025506;
publickey_row[14] = `CIPHERTEXT_WIDTH'd14909164;
publickey_row[15] = `CIPHERTEXT_WIDTH'd4780619;
publickey_row[16] = `CIPHERTEXT_WIDTH'd3882673;
publickey_row[17] = `CIPHERTEXT_WIDTH'd6558100;
publickey_row[18] = `CIPHERTEXT_WIDTH'd8456203;
publickey_row[19] = `CIPHERTEXT_WIDTH'd668712;
publickey_row[20] = `CIPHERTEXT_WIDTH'd3092188;
publickey_row[21] = `CIPHERTEXT_WIDTH'd10008209;
publickey_row[22] = `CIPHERTEXT_WIDTH'd5969800;
publickey_row[23] = `CIPHERTEXT_WIDTH'd15825189;
publickey_row[24] = `CIPHERTEXT_WIDTH'd3177596;
publickey_row[25] = `CIPHERTEXT_WIDTH'd8665256;
publickey_row[26] = `CIPHERTEXT_WIDTH'd10869207;
publickey_row[27] = `CIPHERTEXT_WIDTH'd5879402;
publickey_row[28] = `CIPHERTEXT_WIDTH'd10629024;
publickey_row[29] = `CIPHERTEXT_WIDTH'd12993893;
publickey_row[30] = `CIPHERTEXT_WIDTH'd10527849;
publickey_row[31] = `CIPHERTEXT_WIDTH'd5987403;
publickey_row[32] = `CIPHERTEXT_WIDTH'd1259145;
publickey_row[33] = `CIPHERTEXT_WIDTH'd8933145;
publickey_row[34] = `CIPHERTEXT_WIDTH'd6712985;
publickey_row[35] = `CIPHERTEXT_WIDTH'd6564754;
publickey_row[36] = `CIPHERTEXT_WIDTH'd11111759;
publickey_row[37] = `CIPHERTEXT_WIDTH'd1739197;
publickey_row[38] = `CIPHERTEXT_WIDTH'd12051977;
publickey_row[39] = `CIPHERTEXT_WIDTH'd14233347;
publickey_row[40] = `CIPHERTEXT_WIDTH'd9736314;
publickey_row[41] = `CIPHERTEXT_WIDTH'd539783;
publickey_row[42] = `CIPHERTEXT_WIDTH'd14876748;
publickey_row[43] = `CIPHERTEXT_WIDTH'd4909811;
publickey_row[44] = `CIPHERTEXT_WIDTH'd693722;
publickey_row[45] = `CIPHERTEXT_WIDTH'd15548709;
publickey_row[46] = `CIPHERTEXT_WIDTH'd11589973;
publickey_row[47] = `CIPHERTEXT_WIDTH'd4505500;
publickey_row[48] = `CIPHERTEXT_WIDTH'd8077592;
publickey_row[49] = `CIPHERTEXT_WIDTH'd16770401;
publickey_row[50] = `CIPHERTEXT_WIDTH'd12268114;
publickey_row[51] = `CIPHERTEXT_WIDTH'd13215006;
publickey_row[52] = `CIPHERTEXT_WIDTH'd15409334;
publickey_row[53] = `CIPHERTEXT_WIDTH'd4444515;
publickey_row[54] = `CIPHERTEXT_WIDTH'd1780654;
publickey_row[55] = `CIPHERTEXT_WIDTH'd1631048;
publickey_row[56] = `CIPHERTEXT_WIDTH'd4718345;
publickey_row[57] = `CIPHERTEXT_WIDTH'd7693046;
publickey_row[58] = `CIPHERTEXT_WIDTH'd10657772;
publickey_row[59] = `CIPHERTEXT_WIDTH'd5011322;
publickey_row[60] = `CIPHERTEXT_WIDTH'd11951288;
publickey_row[61] = `CIPHERTEXT_WIDTH'd2630789;
publickey_row[62] = `CIPHERTEXT_WIDTH'd7244619;
publickey_row[63] = `CIPHERTEXT_WIDTH'd15967729;
publickey_row[64] = `CIPHERTEXT_WIDTH'd2698852;
publickey_row[65] = `CIPHERTEXT_WIDTH'd8482367;
publickey_row[66] = `CIPHERTEXT_WIDTH'd11683684;
publickey_row[67] = `CIPHERTEXT_WIDTH'd3960061;
publickey_row[68] = `CIPHERTEXT_WIDTH'd7042834;
publickey_row[69] = `CIPHERTEXT_WIDTH'd15176274;
publickey_row[70] = `CIPHERTEXT_WIDTH'd7780284;
publickey_row[71] = `CIPHERTEXT_WIDTH'd10411182;
publickey_row[72] = `CIPHERTEXT_WIDTH'd9135779;
publickey_row[73] = `CIPHERTEXT_WIDTH'd6836703;
publickey_row[74] = `CIPHERTEXT_WIDTH'd5092500;
publickey_row[75] = `CIPHERTEXT_WIDTH'd3952094;
publickey_row[76] = `CIPHERTEXT_WIDTH'd5323236;
publickey_row[77] = `CIPHERTEXT_WIDTH'd4286690;
publickey_row[78] = `CIPHERTEXT_WIDTH'd7546403;
publickey_row[79] = `CIPHERTEXT_WIDTH'd10412478;
publickey_row[80] = `CIPHERTEXT_WIDTH'd665799;
publickey_row[81] = `CIPHERTEXT_WIDTH'd401483;
publickey_row[82] = `CIPHERTEXT_WIDTH'd9208297;
publickey_row[83] = `CIPHERTEXT_WIDTH'd3904951;
publickey_row[84] = `CIPHERTEXT_WIDTH'd13234387;
publickey_row[85] = `CIPHERTEXT_WIDTH'd550696;
publickey_row[86] = `CIPHERTEXT_WIDTH'd4290481;
publickey_row[87] = `CIPHERTEXT_WIDTH'd3175666;
publickey_row[88] = `CIPHERTEXT_WIDTH'd8484667;
publickey_row[89] = `CIPHERTEXT_WIDTH'd7883862;
publickey_row[90] = `CIPHERTEXT_WIDTH'd1589085;
publickey_row[91] = `CIPHERTEXT_WIDTH'd7060580;
publickey_row[92] = `CIPHERTEXT_WIDTH'd8726748;
publickey_row[93] = `CIPHERTEXT_WIDTH'd9876197;
publickey_row[94] = `CIPHERTEXT_WIDTH'd2597148;
publickey_row[95] = `CIPHERTEXT_WIDTH'd15022288;
publickey_row[96] = `CIPHERTEXT_WIDTH'd15729402;
publickey_row[97] = `CIPHERTEXT_WIDTH'd6300668;
publickey_row[98] = `CIPHERTEXT_WIDTH'd16424650;
publickey_row[99] = `CIPHERTEXT_WIDTH'd4858260;
publickey_row[100] = `CIPHERTEXT_WIDTH'd1982422;
publickey_row[101] = `CIPHERTEXT_WIDTH'd13516035;
publickey_row[102] = `CIPHERTEXT_WIDTH'd11391813;
publickey_row[103] = `CIPHERTEXT_WIDTH'd1872077;
publickey_row[104] = `CIPHERTEXT_WIDTH'd599489;
publickey_row[105] = `CIPHERTEXT_WIDTH'd2341157;
publickey_row[106] = `CIPHERTEXT_WIDTH'd14367642;
publickey_row[107] = `CIPHERTEXT_WIDTH'd428689;
publickey_row[108] = `CIPHERTEXT_WIDTH'd9124702;
publickey_row[109] = `CIPHERTEXT_WIDTH'd4723140;
publickey_row[110] = `CIPHERTEXT_WIDTH'd12273992;
publickey_row[111] = `CIPHERTEXT_WIDTH'd9898216;
publickey_row[112] = `CIPHERTEXT_WIDTH'd10986045;
publickey_row[113] = `CIPHERTEXT_WIDTH'd16079394;
publickey_row[114] = `CIPHERTEXT_WIDTH'd16704336;
publickey_row[115] = `CIPHERTEXT_WIDTH'd13238507;
publickey_row[116] = `CIPHERTEXT_WIDTH'd6044805;
publickey_row[117] = `CIPHERTEXT_WIDTH'd14806709;
publickey_row[118] = `CIPHERTEXT_WIDTH'd6871162;
publickey_row[119] = `CIPHERTEXT_WIDTH'd1640304;
publickey_row[120] = `CIPHERTEXT_WIDTH'd10486142;
publickey_row[121] = `CIPHERTEXT_WIDTH'd8429530;
publickey_row[122] = `CIPHERTEXT_WIDTH'd5360723;
publickey_row[123] = `CIPHERTEXT_WIDTH'd4540327;
publickey_row[124] = `CIPHERTEXT_WIDTH'd10003021;
publickey_row[125] = `CIPHERTEXT_WIDTH'd6523452;
publickey_row[126] = `CIPHERTEXT_WIDTH'd13420732;
publickey_row[127] = `CIPHERTEXT_WIDTH'd12223978;
publickey_row[128] = `CIPHERTEXT_WIDTH'd14401370;
publickey_row[129] = `CIPHERTEXT_WIDTH'd6616173;
publickey_row[130] = `CIPHERTEXT_WIDTH'd2476906;
publickey_row[131] = `CIPHERTEXT_WIDTH'd12934287;
publickey_row[132] = `CIPHERTEXT_WIDTH'd11196015;
publickey_row[133] = `CIPHERTEXT_WIDTH'd4894122;
publickey_row[134] = `CIPHERTEXT_WIDTH'd3532491;
publickey_row[135] = `CIPHERTEXT_WIDTH'd14255436;
publickey_row[136] = `CIPHERTEXT_WIDTH'd4545449;
publickey_row[137] = `CIPHERTEXT_WIDTH'd16509037;
publickey_row[138] = `CIPHERTEXT_WIDTH'd15939970;
publickey_row[139] = `CIPHERTEXT_WIDTH'd6630782;
publickey_row[140] = `CIPHERTEXT_WIDTH'd5446686;
publickey_row[141] = `CIPHERTEXT_WIDTH'd9062563;
publickey_row[142] = `CIPHERTEXT_WIDTH'd11681820;
publickey_row[143] = `CIPHERTEXT_WIDTH'd13335770;
publickey_row[144] = `CIPHERTEXT_WIDTH'd3587980;
publickey_row[145] = `CIPHERTEXT_WIDTH'd7650153;
publickey_row[146] = `CIPHERTEXT_WIDTH'd1717111;
publickey_row[147] = `CIPHERTEXT_WIDTH'd4966488;
publickey_row[148] = `CIPHERTEXT_WIDTH'd8993858;
publickey_row[149] = `CIPHERTEXT_WIDTH'd390172;
publickey_row[150] = `CIPHERTEXT_WIDTH'd9581622;
publickey_row[151] = `CIPHERTEXT_WIDTH'd7381247;
publickey_row[152] = `CIPHERTEXT_WIDTH'd8122888;
publickey_row[153] = `CIPHERTEXT_WIDTH'd8515293;
publickey_row[154] = `CIPHERTEXT_WIDTH'd5295392;
publickey_row[155] = `CIPHERTEXT_WIDTH'd6401072;
publickey_row[156] = `CIPHERTEXT_WIDTH'd2340644;
publickey_row[157] = `CIPHERTEXT_WIDTH'd7104412;
publickey_row[158] = `CIPHERTEXT_WIDTH'd11736728;
publickey_row[159] = `CIPHERTEXT_WIDTH'd7989307;
publickey_row[160] = `CIPHERTEXT_WIDTH'd15515956;
publickey_row[161] = `CIPHERTEXT_WIDTH'd12080773;
publickey_row[162] = `CIPHERTEXT_WIDTH'd10460160;
publickey_row[163] = `CIPHERTEXT_WIDTH'd8223161;
publickey_row[164] = `CIPHERTEXT_WIDTH'd16215350;
publickey_row[165] = `CIPHERTEXT_WIDTH'd14527608;
publickey_row[166] = `CIPHERTEXT_WIDTH'd5382176;
publickey_row[167] = `CIPHERTEXT_WIDTH'd2718538;
publickey_row[168] = `CIPHERTEXT_WIDTH'd2013806;
publickey_row[169] = `CIPHERTEXT_WIDTH'd13838347;
publickey_row[170] = `CIPHERTEXT_WIDTH'd12551524;
publickey_row[171] = `CIPHERTEXT_WIDTH'd9704735;
publickey_row[172] = `CIPHERTEXT_WIDTH'd10948518;
publickey_row[173] = `CIPHERTEXT_WIDTH'd10934120;
publickey_row[174] = `CIPHERTEXT_WIDTH'd10806031;
publickey_row[175] = `CIPHERTEXT_WIDTH'd7921083;
publickey_row[176] = `CIPHERTEXT_WIDTH'd2020774;
publickey_row[177] = `CIPHERTEXT_WIDTH'd2655791;
publickey_row[178] = `CIPHERTEXT_WIDTH'd14977742;
publickey_row[179] = `CIPHERTEXT_WIDTH'd3071369;
publickey_row[180] = `CIPHERTEXT_WIDTH'd4472754;
publickey_row[181] = `CIPHERTEXT_WIDTH'd1226524;
publickey_row[182] = `CIPHERTEXT_WIDTH'd12872850;
publickey_row[183] = `CIPHERTEXT_WIDTH'd206634;
publickey_row[184] = `CIPHERTEXT_WIDTH'd16169471;
publickey_row[185] = `CIPHERTEXT_WIDTH'd2802975;
publickey_row[186] = `CIPHERTEXT_WIDTH'd343957;
publickey_row[187] = `CIPHERTEXT_WIDTH'd15911659;
publickey_row[188] = `CIPHERTEXT_WIDTH'd12031450;
publickey_row[189] = `CIPHERTEXT_WIDTH'd6086630;
publickey_row[190] = `CIPHERTEXT_WIDTH'd3938211;
publickey_row[191] = `CIPHERTEXT_WIDTH'd8893750;
publickey_row[192] = `CIPHERTEXT_WIDTH'd16575883;
publickey_row[193] = `CIPHERTEXT_WIDTH'd11080779;
publickey_row[194] = `CIPHERTEXT_WIDTH'd9041868;
publickey_row[195] = `CIPHERTEXT_WIDTH'd11985321;
publickey_row[196] = `CIPHERTEXT_WIDTH'd16525339;
publickey_row[197] = `CIPHERTEXT_WIDTH'd10779881;
publickey_row[198] = `CIPHERTEXT_WIDTH'd1722864;
publickey_row[199] = `CIPHERTEXT_WIDTH'd9650469;
publickey_row[200] = `CIPHERTEXT_WIDTH'd6346682;
publickey_row[201] = `CIPHERTEXT_WIDTH'd14306249;
publickey_row[202] = `CIPHERTEXT_WIDTH'd8276080;
publickey_row[203] = `CIPHERTEXT_WIDTH'd7376921;
publickey_row[204] = `CIPHERTEXT_WIDTH'd16428230;
publickey_row[205] = `CIPHERTEXT_WIDTH'd2933005;
publickey_row[206] = `CIPHERTEXT_WIDTH'd9961580;
publickey_row[207] = `CIPHERTEXT_WIDTH'd15216328;
publickey_row[208] = `CIPHERTEXT_WIDTH'd9066305;
publickey_row[209] = `CIPHERTEXT_WIDTH'd11966251;
publickey_row[210] = `CIPHERTEXT_WIDTH'd10543672;
publickey_row[211] = `CIPHERTEXT_WIDTH'd830157;
publickey_row[212] = `CIPHERTEXT_WIDTH'd3925906;
publickey_row[213] = `CIPHERTEXT_WIDTH'd5352128;
publickey_row[214] = `CIPHERTEXT_WIDTH'd12101821;
publickey_row[215] = `CIPHERTEXT_WIDTH'd8796607;
publickey_row[216] = `CIPHERTEXT_WIDTH'd7364543;
publickey_row[217] = `CIPHERTEXT_WIDTH'd12984356;
publickey_row[218] = `CIPHERTEXT_WIDTH'd16194162;
publickey_row[219] = `CIPHERTEXT_WIDTH'd9930936;
publickey_row[220] = `CIPHERTEXT_WIDTH'd4804249;
publickey_row[221] = `CIPHERTEXT_WIDTH'd10275208;
publickey_row[222] = `CIPHERTEXT_WIDTH'd6119277;
publickey_row[223] = `CIPHERTEXT_WIDTH'd15975681;
publickey_row[224] = `CIPHERTEXT_WIDTH'd460428;
publickey_row[225] = `CIPHERTEXT_WIDTH'd2296262;
publickey_row[226] = `CIPHERTEXT_WIDTH'd6428129;
publickey_row[227] = `CIPHERTEXT_WIDTH'd11712223;
publickey_row[228] = `CIPHERTEXT_WIDTH'd6399542;
publickey_row[229] = `CIPHERTEXT_WIDTH'd15519375;
publickey_row[230] = `CIPHERTEXT_WIDTH'd5779206;
publickey_row[231] = `CIPHERTEXT_WIDTH'd4610014;
publickey_row[232] = `CIPHERTEXT_WIDTH'd2110802;
publickey_row[233] = `CIPHERTEXT_WIDTH'd12146686;
publickey_row[234] = `CIPHERTEXT_WIDTH'd4194957;
publickey_row[235] = `CIPHERTEXT_WIDTH'd10185867;
publickey_row[236] = `CIPHERTEXT_WIDTH'd12180730;
publickey_row[237] = `CIPHERTEXT_WIDTH'd7860651;
publickey_row[238] = `CIPHERTEXT_WIDTH'd14163609;
publickey_row[239] = `CIPHERTEXT_WIDTH'd2521620;
publickey_row[240] = `CIPHERTEXT_WIDTH'd11863885;
publickey_row[241] = `CIPHERTEXT_WIDTH'd10885514;
publickey_row[242] = `CIPHERTEXT_WIDTH'd4286604;
publickey_row[243] = `CIPHERTEXT_WIDTH'd13901847;
publickey_row[244] = `CIPHERTEXT_WIDTH'd15212398;
publickey_row[245] = `CIPHERTEXT_WIDTH'd3696888;
publickey_row[246] = `CIPHERTEXT_WIDTH'd5116612;
publickey_row[247] = `CIPHERTEXT_WIDTH'd12180923;
publickey_row[248] = `CIPHERTEXT_WIDTH'd10647693;
publickey_row[249] = `CIPHERTEXT_WIDTH'd15444939;
publickey_row[250] = `CIPHERTEXT_WIDTH'd11486975;
publickey_row[251] = `CIPHERTEXT_WIDTH'd1775451;
publickey_row[252] = `CIPHERTEXT_WIDTH'd9995504;
publickey_row[253] = `CIPHERTEXT_WIDTH'd981534;
publickey_row[254] = `CIPHERTEXT_WIDTH'd8441648;
publickey_row[255] = `CIPHERTEXT_WIDTH'd5651076;
publickey_row[256] = `CIPHERTEXT_WIDTH'd11681007;
publickey_row[257] = `CIPHERTEXT_WIDTH'd6071478;
publickey_row[258] = `CIPHERTEXT_WIDTH'd5079858;
publickey_row[259] = `CIPHERTEXT_WIDTH'd15279652;
publickey_row[260] = `CIPHERTEXT_WIDTH'd1479693;
publickey_row[261] = `CIPHERTEXT_WIDTH'd15136727;
publickey_row[262] = `CIPHERTEXT_WIDTH'd12092856;
publickey_row[263] = `CIPHERTEXT_WIDTH'd292021;
publickey_row[264] = `CIPHERTEXT_WIDTH'd13036690;
publickey_row[265] = `CIPHERTEXT_WIDTH'd4023037;
publickey_row[266] = `CIPHERTEXT_WIDTH'd16455610;
publickey_row[267] = `CIPHERTEXT_WIDTH'd2763492;
publickey_row[268] = `CIPHERTEXT_WIDTH'd5794797;
publickey_row[269] = `CIPHERTEXT_WIDTH'd6953642;
publickey_row[270] = `CIPHERTEXT_WIDTH'd14286443;
publickey_row[271] = `CIPHERTEXT_WIDTH'd13931707;
publickey_row[272] = `CIPHERTEXT_WIDTH'd10137969;
publickey_row[273] = `CIPHERTEXT_WIDTH'd6158501;
publickey_row[274] = `CIPHERTEXT_WIDTH'd4810333;
publickey_row[275] = `CIPHERTEXT_WIDTH'd10839460;
publickey_row[276] = `CIPHERTEXT_WIDTH'd10515912;
publickey_row[277] = `CIPHERTEXT_WIDTH'd14548794;
publickey_row[278] = `CIPHERTEXT_WIDTH'd1372513;
publickey_row[279] = `CIPHERTEXT_WIDTH'd11469162;
publickey_row[280] = `CIPHERTEXT_WIDTH'd8729734;
publickey_row[281] = `CIPHERTEXT_WIDTH'd12718943;
publickey_row[282] = `CIPHERTEXT_WIDTH'd5634534;
publickey_row[283] = `CIPHERTEXT_WIDTH'd6311024;
publickey_row[284] = `CIPHERTEXT_WIDTH'd12069437;
publickey_row[285] = `CIPHERTEXT_WIDTH'd13758006;
publickey_row[286] = `CIPHERTEXT_WIDTH'd4156781;
publickey_row[287] = `CIPHERTEXT_WIDTH'd506398;
publickey_row[288] = `CIPHERTEXT_WIDTH'd2623084;
publickey_row[289] = `CIPHERTEXT_WIDTH'd4383965;
publickey_row[290] = `CIPHERTEXT_WIDTH'd8529779;
publickey_row[291] = `CIPHERTEXT_WIDTH'd1559613;
publickey_row[292] = `CIPHERTEXT_WIDTH'd7465933;
publickey_row[293] = `CIPHERTEXT_WIDTH'd4473963;
publickey_row[294] = `CIPHERTEXT_WIDTH'd16085427;
publickey_row[295] = `CIPHERTEXT_WIDTH'd2908614;
publickey_row[296] = `CIPHERTEXT_WIDTH'd13416912;
publickey_row[297] = `CIPHERTEXT_WIDTH'd13273440;
publickey_row[298] = `CIPHERTEXT_WIDTH'd14287662;
publickey_row[299] = `CIPHERTEXT_WIDTH'd10316166;
publickey_row[300] = `CIPHERTEXT_WIDTH'd15161170;
publickey_row[301] = `CIPHERTEXT_WIDTH'd14981131;
publickey_row[302] = `CIPHERTEXT_WIDTH'd2613538;
publickey_row[303] = `CIPHERTEXT_WIDTH'd10613884;
publickey_row[304] = `CIPHERTEXT_WIDTH'd2423527;
publickey_row[305] = `CIPHERTEXT_WIDTH'd11725848;
publickey_row[306] = `CIPHERTEXT_WIDTH'd9103880;
publickey_row[307] = `CIPHERTEXT_WIDTH'd775847;
publickey_row[308] = `CIPHERTEXT_WIDTH'd7311119;
publickey_row[309] = `CIPHERTEXT_WIDTH'd5304193;
publickey_row[310] = `CIPHERTEXT_WIDTH'd12515145;
publickey_row[311] = `CIPHERTEXT_WIDTH'd10266860;
publickey_row[312] = `CIPHERTEXT_WIDTH'd5991591;
publickey_row[313] = `CIPHERTEXT_WIDTH'd4414123;
publickey_row[314] = `CIPHERTEXT_WIDTH'd10451430;
publickey_row[315] = `CIPHERTEXT_WIDTH'd3972226;
publickey_row[316] = `CIPHERTEXT_WIDTH'd10711774;
publickey_row[317] = `CIPHERTEXT_WIDTH'd8056970;
publickey_row[318] = `CIPHERTEXT_WIDTH'd11667206;
publickey_row[319] = `CIPHERTEXT_WIDTH'd13117264;
publickey_row[320] = `CIPHERTEXT_WIDTH'd1658956;
publickey_row[321] = `CIPHERTEXT_WIDTH'd2034976;
publickey_row[322] = `CIPHERTEXT_WIDTH'd12596020;
publickey_row[323] = `CIPHERTEXT_WIDTH'd15664250;
publickey_row[324] = `CIPHERTEXT_WIDTH'd12511461;
publickey_row[325] = `CIPHERTEXT_WIDTH'd4333422;
publickey_row[326] = `CIPHERTEXT_WIDTH'd13471456;
publickey_row[327] = `CIPHERTEXT_WIDTH'd16615098;
publickey_row[328] = `CIPHERTEXT_WIDTH'd264108;
publickey_row[329] = `CIPHERTEXT_WIDTH'd1822032;
publickey_row[330] = `CIPHERTEXT_WIDTH'd10158433;
publickey_row[331] = `CIPHERTEXT_WIDTH'd7321578;
publickey_row[332] = `CIPHERTEXT_WIDTH'd1739769;
publickey_row[333] = `CIPHERTEXT_WIDTH'd12860666;
publickey_row[334] = `CIPHERTEXT_WIDTH'd4539498;
publickey_row[335] = `CIPHERTEXT_WIDTH'd3145358;
publickey_row[336] = `CIPHERTEXT_WIDTH'd5512727;
publickey_row[337] = `CIPHERTEXT_WIDTH'd11669050;
publickey_row[338] = `CIPHERTEXT_WIDTH'd11149823;
publickey_row[339] = `CIPHERTEXT_WIDTH'd7470229;
publickey_row[340] = `CIPHERTEXT_WIDTH'd11598480;
publickey_row[341] = `CIPHERTEXT_WIDTH'd6462320;
publickey_row[342] = `CIPHERTEXT_WIDTH'd12432519;
publickey_row[343] = `CIPHERTEXT_WIDTH'd7024080;
publickey_row[344] = `CIPHERTEXT_WIDTH'd7861084;
publickey_row[345] = `CIPHERTEXT_WIDTH'd14671106;
publickey_row[346] = `CIPHERTEXT_WIDTH'd15341892;
publickey_row[347] = `CIPHERTEXT_WIDTH'd6153096;
publickey_row[348] = `CIPHERTEXT_WIDTH'd16220841;
publickey_row[349] = `CIPHERTEXT_WIDTH'd6846510;
publickey_row[350] = `CIPHERTEXT_WIDTH'd12649304;
publickey_row[351] = `CIPHERTEXT_WIDTH'd4216508;
publickey_row[352] = `CIPHERTEXT_WIDTH'd590769;
publickey_row[353] = `CIPHERTEXT_WIDTH'd13240174;
publickey_row[354] = `CIPHERTEXT_WIDTH'd16083680;
publickey_row[355] = `CIPHERTEXT_WIDTH'd4884102;
publickey_row[356] = `CIPHERTEXT_WIDTH'd6216489;
publickey_row[357] = `CIPHERTEXT_WIDTH'd11339654;
publickey_row[358] = `CIPHERTEXT_WIDTH'd11496255;
publickey_row[359] = `CIPHERTEXT_WIDTH'd6782867;
publickey_row[360] = `CIPHERTEXT_WIDTH'd10289595;
publickey_row[361] = `CIPHERTEXT_WIDTH'd11196147;
publickey_row[362] = `CIPHERTEXT_WIDTH'd5194297;
publickey_row[363] = `CIPHERTEXT_WIDTH'd13613839;
publickey_row[364] = `CIPHERTEXT_WIDTH'd11282105;
publickey_row[365] = `CIPHERTEXT_WIDTH'd14342531;
publickey_row[366] = `CIPHERTEXT_WIDTH'd2865737;
publickey_row[367] = `CIPHERTEXT_WIDTH'd16375219;
publickey_row[368] = `CIPHERTEXT_WIDTH'd8527524;
publickey_row[369] = `CIPHERTEXT_WIDTH'd7117667;
publickey_row[370] = `CIPHERTEXT_WIDTH'd11838431;
publickey_row[371] = `CIPHERTEXT_WIDTH'd5194478;
publickey_row[372] = `CIPHERTEXT_WIDTH'd13222861;
publickey_row[373] = `CIPHERTEXT_WIDTH'd6234059;
publickey_row[374] = `CIPHERTEXT_WIDTH'd9034285;
publickey_row[375] = `CIPHERTEXT_WIDTH'd11044728;
publickey_row[376] = `CIPHERTEXT_WIDTH'd5802168;
publickey_row[377] = `CIPHERTEXT_WIDTH'd8855929;
publickey_row[378] = `CIPHERTEXT_WIDTH'd14317962;
publickey_row[379] = `CIPHERTEXT_WIDTH'd12231546;
publickey_row[380] = `CIPHERTEXT_WIDTH'd12064375;
publickey_row[381] = `CIPHERTEXT_WIDTH'd12493375;
publickey_row[382] = `CIPHERTEXT_WIDTH'd7910344;
publickey_row[383] = `CIPHERTEXT_WIDTH'd11510397;
publickey_row[384] = `CIPHERTEXT_WIDTH'd3631739;
publickey_row[385] = `CIPHERTEXT_WIDTH'd12606761;
publickey_row[386] = `CIPHERTEXT_WIDTH'd10726673;
publickey_row[387] = `CIPHERTEXT_WIDTH'd15435532;
publickey_row[388] = `CIPHERTEXT_WIDTH'd11123706;
publickey_row[389] = `CIPHERTEXT_WIDTH'd16537536;
publickey_row[390] = `CIPHERTEXT_WIDTH'd12469602;
publickey_row[391] = `CIPHERTEXT_WIDTH'd3010808;
publickey_row[392] = `CIPHERTEXT_WIDTH'd5182098;
publickey_row[393] = `CIPHERTEXT_WIDTH'd11068622;
publickey_row[394] = `CIPHERTEXT_WIDTH'd6338665;
publickey_row[395] = `CIPHERTEXT_WIDTH'd3828927;
publickey_row[396] = `CIPHERTEXT_WIDTH'd6846790;
publickey_row[397] = `CIPHERTEXT_WIDTH'd1898815;
publickey_row[398] = `CIPHERTEXT_WIDTH'd11890537;
publickey_row[399] = `CIPHERTEXT_WIDTH'd10895854;
publickey_row[400] = `CIPHERTEXT_WIDTH'd12310682;
publickey_row[401] = `CIPHERTEXT_WIDTH'd3007458;
publickey_row[402] = `CIPHERTEXT_WIDTH'd15697212;
publickey_row[403] = `CIPHERTEXT_WIDTH'd11295215;
publickey_row[404] = `CIPHERTEXT_WIDTH'd13651966;
publickey_row[405] = `CIPHERTEXT_WIDTH'd4968476;
publickey_row[406] = `CIPHERTEXT_WIDTH'd10532548;
publickey_row[407] = `CIPHERTEXT_WIDTH'd13891661;
publickey_row[408] = `CIPHERTEXT_WIDTH'd11514806;
publickey_row[409] = `CIPHERTEXT_WIDTH'd16166319;
publickey_row[410] = `CIPHERTEXT_WIDTH'd51737;
publickey_row[411] = `CIPHERTEXT_WIDTH'd11946565;
publickey_row[412] = `CIPHERTEXT_WIDTH'd12114329;
publickey_row[413] = `CIPHERTEXT_WIDTH'd2180529;
publickey_row[414] = `CIPHERTEXT_WIDTH'd11627830;
publickey_row[415] = `CIPHERTEXT_WIDTH'd1343163;
publickey_row[416] = `CIPHERTEXT_WIDTH'd11526150;
publickey_row[417] = `CIPHERTEXT_WIDTH'd12029382;
publickey_row[418] = `CIPHERTEXT_WIDTH'd14689717;
publickey_row[419] = `CIPHERTEXT_WIDTH'd13138288;
publickey_row[420] = `CIPHERTEXT_WIDTH'd3414236;
publickey_row[421] = `CIPHERTEXT_WIDTH'd4576688;
publickey_row[422] = `CIPHERTEXT_WIDTH'd6478690;
publickey_row[423] = `CIPHERTEXT_WIDTH'd1320622;
publickey_row[424] = `CIPHERTEXT_WIDTH'd7655006;
publickey_row[425] = `CIPHERTEXT_WIDTH'd8455609;
publickey_row[426] = `CIPHERTEXT_WIDTH'd7186756;
publickey_row[427] = `CIPHERTEXT_WIDTH'd4084998;
publickey_row[428] = `CIPHERTEXT_WIDTH'd8680426;
publickey_row[429] = `CIPHERTEXT_WIDTH'd8810168;
publickey_row[430] = `CIPHERTEXT_WIDTH'd10960225;
publickey_row[431] = `CIPHERTEXT_WIDTH'd7810277;
publickey_row[432] = `CIPHERTEXT_WIDTH'd11850484;
publickey_row[433] = `CIPHERTEXT_WIDTH'd16450357;
publickey_row[434] = `CIPHERTEXT_WIDTH'd5874573;
publickey_row[435] = `CIPHERTEXT_WIDTH'd5174554;
publickey_row[436] = `CIPHERTEXT_WIDTH'd12773526;
publickey_row[437] = `CIPHERTEXT_WIDTH'd11447391;
publickey_row[438] = `CIPHERTEXT_WIDTH'd2905343;
publickey_row[439] = `CIPHERTEXT_WIDTH'd15878695;
publickey_row[440] = `CIPHERTEXT_WIDTH'd3656883;
publickey_row[441] = `CIPHERTEXT_WIDTH'd5258049;
publickey_row[442] = `CIPHERTEXT_WIDTH'd8554470;
publickey_row[443] = `CIPHERTEXT_WIDTH'd2699060;
publickey_row[444] = `CIPHERTEXT_WIDTH'd6379958;
publickey_row[445] = `CIPHERTEXT_WIDTH'd1195443;
publickey_row[446] = `CIPHERTEXT_WIDTH'd14086088;
publickey_row[447] = `CIPHERTEXT_WIDTH'd11351843;
publickey_row[448] = `CIPHERTEXT_WIDTH'd8671360;
publickey_row[449] = `CIPHERTEXT_WIDTH'd5167691;
publickey_row[450] = `CIPHERTEXT_WIDTH'd1346588;
publickey_row[451] = `CIPHERTEXT_WIDTH'd815254;
publickey_row[452] = `CIPHERTEXT_WIDTH'd3627117;
publickey_row[453] = `CIPHERTEXT_WIDTH'd4311050;
publickey_row[454] = `CIPHERTEXT_WIDTH'd3242342;
publickey_row[455] = `CIPHERTEXT_WIDTH'd12189088;
publickey_row[456] = `CIPHERTEXT_WIDTH'd15939262;
publickey_row[457] = `CIPHERTEXT_WIDTH'd14333713;
publickey_row[458] = `CIPHERTEXT_WIDTH'd6200461;
publickey_row[459] = `CIPHERTEXT_WIDTH'd8630235;
publickey_row[460] = `CIPHERTEXT_WIDTH'd13067448;
publickey_row[461] = `CIPHERTEXT_WIDTH'd12754734;
publickey_row[462] = `CIPHERTEXT_WIDTH'd2375560;
publickey_row[463] = `CIPHERTEXT_WIDTH'd10009108;
publickey_row[464] = `CIPHERTEXT_WIDTH'd11043139;
publickey_row[465] = `CIPHERTEXT_WIDTH'd3744652;
publickey_row[466] = `CIPHERTEXT_WIDTH'd6151622;
publickey_row[467] = `CIPHERTEXT_WIDTH'd11926411;
publickey_row[468] = `CIPHERTEXT_WIDTH'd9496903;
publickey_row[469] = `CIPHERTEXT_WIDTH'd2415893;
publickey_row[470] = `CIPHERTEXT_WIDTH'd3961494;
publickey_row[471] = `CIPHERTEXT_WIDTH'd9672708;
publickey_row[472] = `CIPHERTEXT_WIDTH'd9461367;
publickey_row[473] = `CIPHERTEXT_WIDTH'd8299153;
publickey_row[474] = `CIPHERTEXT_WIDTH'd5676173;
publickey_row[475] = `CIPHERTEXT_WIDTH'd3409518;
publickey_row[476] = `CIPHERTEXT_WIDTH'd4181144;
publickey_row[477] = `CIPHERTEXT_WIDTH'd7284157;
publickey_row[478] = `CIPHERTEXT_WIDTH'd15149121;
publickey_row[479] = `CIPHERTEXT_WIDTH'd7618866;
publickey_row[480] = `CIPHERTEXT_WIDTH'd16505156;
publickey_row[481] = `CIPHERTEXT_WIDTH'd5884859;
publickey_row[482] = `CIPHERTEXT_WIDTH'd67926;
publickey_row[483] = `CIPHERTEXT_WIDTH'd14747928;
publickey_row[484] = `CIPHERTEXT_WIDTH'd9309757;
publickey_row[485] = `CIPHERTEXT_WIDTH'd9282705;
publickey_row[486] = `CIPHERTEXT_WIDTH'd6998316;
publickey_row[487] = `CIPHERTEXT_WIDTH'd9962602;
publickey_row[488] = `CIPHERTEXT_WIDTH'd15458533;
publickey_row[489] = `CIPHERTEXT_WIDTH'd10032893;
publickey_row[490] = `CIPHERTEXT_WIDTH'd2232395;
publickey_row[491] = `CIPHERTEXT_WIDTH'd12929286;
publickey_row[492] = `CIPHERTEXT_WIDTH'd2744855;
publickey_row[493] = `CIPHERTEXT_WIDTH'd2068248;
publickey_row[494] = `CIPHERTEXT_WIDTH'd8874962;
publickey_row[495] = `CIPHERTEXT_WIDTH'd3435366;
publickey_row[496] = `CIPHERTEXT_WIDTH'd11563490;
publickey_row[497] = `CIPHERTEXT_WIDTH'd10884959;
publickey_row[498] = `CIPHERTEXT_WIDTH'd13001051;
publickey_row[499] = `CIPHERTEXT_WIDTH'd3909542;
publickey_row[500] = `CIPHERTEXT_WIDTH'd2042022;
publickey_row[501] = `CIPHERTEXT_WIDTH'd3819500;
publickey_row[502] = `CIPHERTEXT_WIDTH'd11760955;
publickey_row[503] = `CIPHERTEXT_WIDTH'd16313520;
publickey_row[504] = `CIPHERTEXT_WIDTH'd12311526;
publickey_row[505] = `CIPHERTEXT_WIDTH'd3246859;
publickey_row[506] = `CIPHERTEXT_WIDTH'd1346284;
publickey_row[507] = `CIPHERTEXT_WIDTH'd12629248;
publickey_row[508] = `CIPHERTEXT_WIDTH'd8695237;
publickey_row[509] = `CIPHERTEXT_WIDTH'd7584833;
publickey_row[510] = `CIPHERTEXT_WIDTH'd8256480;
publickey_row[511] = `CIPHERTEXT_WIDTH'd14126582;
publickey_row[512] = `CIPHERTEXT_WIDTH'd881716;
publickey_row[513] = `CIPHERTEXT_WIDTH'd9224668;
publickey_row[514] = `CIPHERTEXT_WIDTH'd6109401;
publickey_row[515] = `CIPHERTEXT_WIDTH'd2471639;
publickey_row[516] = `CIPHERTEXT_WIDTH'd12014284;
publickey_row[517] = `CIPHERTEXT_WIDTH'd10104158;
publickey_row[518] = `CIPHERTEXT_WIDTH'd2697691;
publickey_row[519] = `CIPHERTEXT_WIDTH'd11070015;
publickey_row[520] = `CIPHERTEXT_WIDTH'd8077085;
publickey_row[521] = `CIPHERTEXT_WIDTH'd10079540;
publickey_row[522] = `CIPHERTEXT_WIDTH'd12612501;
publickey_row[523] = `CIPHERTEXT_WIDTH'd13337554;
publickey_row[524] = `CIPHERTEXT_WIDTH'd2817971;
publickey_row[525] = `CIPHERTEXT_WIDTH'd10401742;
publickey_row[526] = `CIPHERTEXT_WIDTH'd5671384;
publickey_row[527] = `CIPHERTEXT_WIDTH'd10972057;
publickey_row[528] = `CIPHERTEXT_WIDTH'd9959607;
publickey_row[529] = `CIPHERTEXT_WIDTH'd8530112;
publickey_row[530] = `CIPHERTEXT_WIDTH'd8999948;
publickey_row[531] = `CIPHERTEXT_WIDTH'd1070163;
publickey_row[532] = `CIPHERTEXT_WIDTH'd11251782;
publickey_row[533] = `CIPHERTEXT_WIDTH'd3642641;
publickey_row[534] = `CIPHERTEXT_WIDTH'd16220660;
publickey_row[535] = `CIPHERTEXT_WIDTH'd7344836;
publickey_row[536] = `CIPHERTEXT_WIDTH'd13199347;
publickey_row[537] = `CIPHERTEXT_WIDTH'd9530128;
publickey_row[538] = `CIPHERTEXT_WIDTH'd5479717;
publickey_row[539] = `CIPHERTEXT_WIDTH'd8100317;
publickey_row[540] = `CIPHERTEXT_WIDTH'd11973396;
publickey_row[541] = `CIPHERTEXT_WIDTH'd6480735;
publickey_row[542] = `CIPHERTEXT_WIDTH'd11898643;
publickey_row[543] = `CIPHERTEXT_WIDTH'd2455972;
publickey_row[544] = `CIPHERTEXT_WIDTH'd10202347;
publickey_row[545] = `CIPHERTEXT_WIDTH'd2188909;
publickey_row[546] = `CIPHERTEXT_WIDTH'd11282467;
publickey_row[547] = `CIPHERTEXT_WIDTH'd1550601;
publickey_row[548] = `CIPHERTEXT_WIDTH'd4160138;
publickey_row[549] = `CIPHERTEXT_WIDTH'd1516087;
publickey_row[550] = `CIPHERTEXT_WIDTH'd8907051;
publickey_row[551] = `CIPHERTEXT_WIDTH'd4340628;
publickey_row[552] = `CIPHERTEXT_WIDTH'd12879787;
publickey_row[553] = `CIPHERTEXT_WIDTH'd15140697;
publickey_row[554] = `CIPHERTEXT_WIDTH'd14171755;
publickey_row[555] = `CIPHERTEXT_WIDTH'd7396533;
publickey_row[556] = `CIPHERTEXT_WIDTH'd12179473;
publickey_row[557] = `CIPHERTEXT_WIDTH'd11828494;
publickey_row[558] = `CIPHERTEXT_WIDTH'd5922778;
publickey_row[559] = `CIPHERTEXT_WIDTH'd11629343;
publickey_row[560] = `CIPHERTEXT_WIDTH'd11659175;
publickey_row[561] = `CIPHERTEXT_WIDTH'd13330253;
publickey_row[562] = `CIPHERTEXT_WIDTH'd5706644;
publickey_row[563] = `CIPHERTEXT_WIDTH'd8539515;
publickey_row[564] = `CIPHERTEXT_WIDTH'd8172371;
publickey_row[565] = `CIPHERTEXT_WIDTH'd6639695;
publickey_row[566] = `CIPHERTEXT_WIDTH'd1482822;
publickey_row[567] = `CIPHERTEXT_WIDTH'd3183977;
publickey_row[568] = `CIPHERTEXT_WIDTH'd3852985;
publickey_row[569] = `CIPHERTEXT_WIDTH'd15474272;
publickey_row[570] = `CIPHERTEXT_WIDTH'd11780848;
publickey_row[571] = `CIPHERTEXT_WIDTH'd14038969;
publickey_row[572] = `CIPHERTEXT_WIDTH'd1610864;
publickey_row[573] = `CIPHERTEXT_WIDTH'd14891992;
publickey_row[574] = `CIPHERTEXT_WIDTH'd13956860;
publickey_row[575] = `CIPHERTEXT_WIDTH'd750620;
publickey_row[576] = `CIPHERTEXT_WIDTH'd4473387;
publickey_row[577] = `CIPHERTEXT_WIDTH'd16050117;
publickey_row[578] = `CIPHERTEXT_WIDTH'd8502778;
publickey_row[579] = `CIPHERTEXT_WIDTH'd9518515;
publickey_row[580] = `CIPHERTEXT_WIDTH'd649483;
publickey_row[581] = `CIPHERTEXT_WIDTH'd8980912;
publickey_row[582] = `CIPHERTEXT_WIDTH'd15321173;
publickey_row[583] = `CIPHERTEXT_WIDTH'd5244230;
publickey_row[584] = `CIPHERTEXT_WIDTH'd8178082;
publickey_row[585] = `CIPHERTEXT_WIDTH'd1390411;
publickey_row[586] = `CIPHERTEXT_WIDTH'd1266834;
publickey_row[587] = `CIPHERTEXT_WIDTH'd2644984;
publickey_row[588] = `CIPHERTEXT_WIDTH'd11944393;
publickey_row[589] = `CIPHERTEXT_WIDTH'd3729266;
publickey_row[590] = `CIPHERTEXT_WIDTH'd2702358;
publickey_row[591] = `CIPHERTEXT_WIDTH'd5314375;
publickey_row[592] = `CIPHERTEXT_WIDTH'd9624038;
publickey_row[593] = `CIPHERTEXT_WIDTH'd8178253;
publickey_row[594] = `CIPHERTEXT_WIDTH'd3042284;
publickey_row[595] = `CIPHERTEXT_WIDTH'd16230401;
publickey_row[596] = `CIPHERTEXT_WIDTH'd15162274;
publickey_row[597] = `CIPHERTEXT_WIDTH'd7911494;
publickey_row[598] = `CIPHERTEXT_WIDTH'd3714258;
publickey_row[599] = `CIPHERTEXT_WIDTH'd14651586;
publickey_row[600] = `CIPHERTEXT_WIDTH'd4235909;
publickey_row[601] = `CIPHERTEXT_WIDTH'd4296147;
publickey_row[602] = `CIPHERTEXT_WIDTH'd1354820;
publickey_row[603] = `CIPHERTEXT_WIDTH'd728314;
publickey_row[604] = `CIPHERTEXT_WIDTH'd4831335;
publickey_row[605] = `CIPHERTEXT_WIDTH'd71692;
publickey_row[606] = `CIPHERTEXT_WIDTH'd11221416;
publickey_row[607] = `CIPHERTEXT_WIDTH'd10067252;
publickey_row[608] = `CIPHERTEXT_WIDTH'd5981130;
publickey_row[609] = `CIPHERTEXT_WIDTH'd9641693;
publickey_row[610] = `CIPHERTEXT_WIDTH'd13115526;
publickey_row[611] = `CIPHERTEXT_WIDTH'd11152703;
publickey_row[612] = `CIPHERTEXT_WIDTH'd8426223;
publickey_row[613] = `CIPHERTEXT_WIDTH'd3007931;
publickey_row[614] = `CIPHERTEXT_WIDTH'd7653999;
publickey_row[615] = `CIPHERTEXT_WIDTH'd5109266;
publickey_row[616] = `CIPHERTEXT_WIDTH'd1341150;
publickey_row[617] = `CIPHERTEXT_WIDTH'd4659860;
publickey_row[618] = `CIPHERTEXT_WIDTH'd1924383;
publickey_row[619] = `CIPHERTEXT_WIDTH'd9667426;
publickey_row[620] = `CIPHERTEXT_WIDTH'd14191121;
publickey_row[621] = `CIPHERTEXT_WIDTH'd16320036;
publickey_row[622] = `CIPHERTEXT_WIDTH'd14889958;
publickey_row[623] = `CIPHERTEXT_WIDTH'd12700858;
publickey_row[624] = `CIPHERTEXT_WIDTH'd12433829;
publickey_row[625] = `CIPHERTEXT_WIDTH'd1655451;
publickey_row[626] = `CIPHERTEXT_WIDTH'd10466724;
publickey_row[627] = `CIPHERTEXT_WIDTH'd5459828;
publickey_row[628] = `CIPHERTEXT_WIDTH'd9897867;
publickey_row[629] = `CIPHERTEXT_WIDTH'd13198600;
publickey_row[630] = `CIPHERTEXT_WIDTH'd8132042;
publickey_row[631] = `CIPHERTEXT_WIDTH'd3523174;
publickey_row[632] = `CIPHERTEXT_WIDTH'd10570146;
publickey_row[633] = `CIPHERTEXT_WIDTH'd3710928;
publickey_row[634] = `CIPHERTEXT_WIDTH'd15579840;
publickey_row[635] = `CIPHERTEXT_WIDTH'd7140781;
publickey_row[636] = `CIPHERTEXT_WIDTH'd12118582;
publickey_row[637] = `CIPHERTEXT_WIDTH'd16609278;
publickey_row[638] = `CIPHERTEXT_WIDTH'd15335790;
publickey_row[639] = `CIPHERTEXT_WIDTH'd16708150;
publickey_row[640] = `CIPHERTEXT_WIDTH'd15164357;
publickey_row[641] = `CIPHERTEXT_WIDTH'd6100390;
publickey_row[642] = `CIPHERTEXT_WIDTH'd9013174;
publickey_row[643] = `CIPHERTEXT_WIDTH'd6547078;
publickey_row[644] = `CIPHERTEXT_WIDTH'd12566327;
publickey_row[645] = `CIPHERTEXT_WIDTH'd14609734;
publickey_row[646] = `CIPHERTEXT_WIDTH'd970033;
publickey_row[647] = `CIPHERTEXT_WIDTH'd11729700;
publickey_row[648] = `CIPHERTEXT_WIDTH'd10993801;
publickey_row[649] = `CIPHERTEXT_WIDTH'd14737157;
publickey_row[650] = `CIPHERTEXT_WIDTH'd3233682;
publickey_row[651] = `CIPHERTEXT_WIDTH'd9317640;
publickey_row[652] = `CIPHERTEXT_WIDTH'd2330264;
publickey_row[653] = `CIPHERTEXT_WIDTH'd16279450;
publickey_row[654] = `CIPHERTEXT_WIDTH'd11248865;
publickey_row[655] = `CIPHERTEXT_WIDTH'd3573950;
publickey_row[656] = `CIPHERTEXT_WIDTH'd15877601;
publickey_row[657] = `CIPHERTEXT_WIDTH'd16456848;
publickey_row[658] = `CIPHERTEXT_WIDTH'd5944529;
publickey_row[659] = `CIPHERTEXT_WIDTH'd4379520;
publickey_row[660] = `CIPHERTEXT_WIDTH'd13357769;
publickey_row[661] = `CIPHERTEXT_WIDTH'd11190556;
publickey_row[662] = `CIPHERTEXT_WIDTH'd14662814;
publickey_row[663] = `CIPHERTEXT_WIDTH'd8828945;
publickey_row[664] = `CIPHERTEXT_WIDTH'd9915594;
publickey_row[665] = `CIPHERTEXT_WIDTH'd5588601;
publickey_row[666] = `CIPHERTEXT_WIDTH'd15477130;
publickey_row[667] = `CIPHERTEXT_WIDTH'd14928832;
publickey_row[668] = `CIPHERTEXT_WIDTH'd8314649;
publickey_row[669] = `CIPHERTEXT_WIDTH'd5055438;
publickey_row[670] = `CIPHERTEXT_WIDTH'd5044119;
publickey_row[671] = `CIPHERTEXT_WIDTH'd8885145;
publickey_row[672] = `CIPHERTEXT_WIDTH'd612126;
publickey_row[673] = `CIPHERTEXT_WIDTH'd11238052;
publickey_row[674] = `CIPHERTEXT_WIDTH'd6032793;
publickey_row[675] = `CIPHERTEXT_WIDTH'd1314580;
publickey_row[676] = `CIPHERTEXT_WIDTH'd9802573;
publickey_row[677] = `CIPHERTEXT_WIDTH'd14354175;
publickey_row[678] = `CIPHERTEXT_WIDTH'd6664375;
publickey_row[679] = `CIPHERTEXT_WIDTH'd7501992;
publickey_row[680] = `CIPHERTEXT_WIDTH'd13195901;
publickey_row[681] = `CIPHERTEXT_WIDTH'd7440534;
publickey_row[682] = `CIPHERTEXT_WIDTH'd12893927;
publickey_row[683] = `CIPHERTEXT_WIDTH'd4039616;
publickey_row[684] = `CIPHERTEXT_WIDTH'd16404;
publickey_row[685] = `CIPHERTEXT_WIDTH'd8405912;
publickey_row[686] = `CIPHERTEXT_WIDTH'd5857404;
publickey_row[687] = `CIPHERTEXT_WIDTH'd10079524;
publickey_row[688] = `CIPHERTEXT_WIDTH'd12178128;
publickey_row[689] = `CIPHERTEXT_WIDTH'd9783811;
publickey_row[690] = `CIPHERTEXT_WIDTH'd1718230;
publickey_row[691] = `CIPHERTEXT_WIDTH'd6824047;
publickey_row[692] = `CIPHERTEXT_WIDTH'd3359948;
publickey_row[693] = `CIPHERTEXT_WIDTH'd13940581;
publickey_row[694] = `CIPHERTEXT_WIDTH'd3809786;
publickey_row[695] = `CIPHERTEXT_WIDTH'd4799254;
publickey_row[696] = `CIPHERTEXT_WIDTH'd11672182;
publickey_row[697] = `CIPHERTEXT_WIDTH'd3760456;
publickey_row[698] = `CIPHERTEXT_WIDTH'd16557861;
publickey_row[699] = `CIPHERTEXT_WIDTH'd9564624;
publickey_row[700] = `CIPHERTEXT_WIDTH'd4223456;
publickey_row[701] = `CIPHERTEXT_WIDTH'd761501;
publickey_row[702] = `CIPHERTEXT_WIDTH'd11484995;
publickey_row[703] = `CIPHERTEXT_WIDTH'd7445694;
publickey_row[704] = `CIPHERTEXT_WIDTH'd15456923;
publickey_row[705] = `CIPHERTEXT_WIDTH'd11843762;
publickey_row[706] = `CIPHERTEXT_WIDTH'd5659375;
publickey_row[707] = `CIPHERTEXT_WIDTH'd5318177;
publickey_row[708] = `CIPHERTEXT_WIDTH'd11820261;
publickey_row[709] = `CIPHERTEXT_WIDTH'd8352470;
publickey_row[710] = `CIPHERTEXT_WIDTH'd8489702;
publickey_row[711] = `CIPHERTEXT_WIDTH'd14521837;
publickey_row[712] = `CIPHERTEXT_WIDTH'd9055300;
publickey_row[713] = `CIPHERTEXT_WIDTH'd12813630;
publickey_row[714] = `CIPHERTEXT_WIDTH'd13093176;
publickey_row[715] = `CIPHERTEXT_WIDTH'd8070955;
publickey_row[716] = `CIPHERTEXT_WIDTH'd9557631;
publickey_row[717] = `CIPHERTEXT_WIDTH'd3422815;
publickey_row[718] = `CIPHERTEXT_WIDTH'd9473782;
publickey_row[719] = `CIPHERTEXT_WIDTH'd215756;
publickey_row[720] = `CIPHERTEXT_WIDTH'd784906;
publickey_row[721] = `CIPHERTEXT_WIDTH'd8372002;
publickey_row[722] = `CIPHERTEXT_WIDTH'd14793871;
publickey_row[723] = `CIPHERTEXT_WIDTH'd15136473;
publickey_row[724] = `CIPHERTEXT_WIDTH'd2980218;
publickey_row[725] = `CIPHERTEXT_WIDTH'd3459615;
publickey_row[726] = `CIPHERTEXT_WIDTH'd13702487;
publickey_row[727] = `CIPHERTEXT_WIDTH'd9532189;
publickey_row[728] = `CIPHERTEXT_WIDTH'd8611090;
publickey_row[729] = `CIPHERTEXT_WIDTH'd8123742;
publickey_row[730] = `CIPHERTEXT_WIDTH'd6698501;
publickey_row[731] = `CIPHERTEXT_WIDTH'd13969044;
publickey_row[732] = `CIPHERTEXT_WIDTH'd3907622;
publickey_row[733] = `CIPHERTEXT_WIDTH'd3815483;
publickey_row[734] = `CIPHERTEXT_WIDTH'd894238;
publickey_row[735] = `CIPHERTEXT_WIDTH'd15693992;
publickey_row[736] = `CIPHERTEXT_WIDTH'd4890398;
publickey_row[737] = `CIPHERTEXT_WIDTH'd7604905;
publickey_row[738] = `CIPHERTEXT_WIDTH'd6367778;
publickey_row[739] = `CIPHERTEXT_WIDTH'd15151407;
publickey_row[740] = `CIPHERTEXT_WIDTH'd3044423;
publickey_row[741] = `CIPHERTEXT_WIDTH'd7287911;
publickey_row[742] = `CIPHERTEXT_WIDTH'd13472164;
publickey_row[743] = `CIPHERTEXT_WIDTH'd10420208;
publickey_row[744] = `CIPHERTEXT_WIDTH'd5123067;
publickey_row[745] = `CIPHERTEXT_WIDTH'd7151160;
publickey_row[746] = `CIPHERTEXT_WIDTH'd4325807;
publickey_row[747] = `CIPHERTEXT_WIDTH'd3464221;
publickey_row[748] = `CIPHERTEXT_WIDTH'd13951721;
publickey_row[749] = `CIPHERTEXT_WIDTH'd15901366;
publickey_row[750] = `CIPHERTEXT_WIDTH'd10592080;
publickey_row[751] = `CIPHERTEXT_WIDTH'd14106985;
publickey_row[752] = `CIPHERTEXT_WIDTH'd15688457;
publickey_row[753] = `CIPHERTEXT_WIDTH'd8731677;
publickey_row[754] = `CIPHERTEXT_WIDTH'd8831742;
publickey_row[755] = `CIPHERTEXT_WIDTH'd6610913;
publickey_row[756] = `CIPHERTEXT_WIDTH'd16092274;
publickey_row[757] = `CIPHERTEXT_WIDTH'd14954003;
publickey_row[758] = `CIPHERTEXT_WIDTH'd10248219;
publickey_row[759] = `CIPHERTEXT_WIDTH'd10906240;
publickey_row[760] = `CIPHERTEXT_WIDTH'd16068454;
publickey_row[761] = `CIPHERTEXT_WIDTH'd13140715;
publickey_row[762] = `CIPHERTEXT_WIDTH'd2692092;
publickey_row[763] = `CIPHERTEXT_WIDTH'd16607828;
publickey_row[764] = `CIPHERTEXT_WIDTH'd14960539;
publickey_row[765] = `CIPHERTEXT_WIDTH'd11744638;
publickey_row[766] = `CIPHERTEXT_WIDTH'd1028207;
publickey_row[767] = `CIPHERTEXT_WIDTH'd7670772;
publickey_row[768] = `CIPHERTEXT_WIDTH'd2105566;
publickey_row[769] = `CIPHERTEXT_WIDTH'd9299082;
publickey_row[770] = `CIPHERTEXT_WIDTH'd16173451;
publickey_row[771] = `CIPHERTEXT_WIDTH'd9398708;
publickey_row[772] = `CIPHERTEXT_WIDTH'd11399145;
publickey_row[773] = `CIPHERTEXT_WIDTH'd7317372;
publickey_row[774] = `CIPHERTEXT_WIDTH'd14196445;
publickey_row[775] = `CIPHERTEXT_WIDTH'd3755431;
publickey_row[776] = `CIPHERTEXT_WIDTH'd4436836;
publickey_row[777] = `CIPHERTEXT_WIDTH'd4699045;
publickey_row[778] = `CIPHERTEXT_WIDTH'd9341744;
publickey_row[779] = `CIPHERTEXT_WIDTH'd9099197;
publickey_row[780] = `CIPHERTEXT_WIDTH'd16139639;
publickey_row[781] = `CIPHERTEXT_WIDTH'd10724738;
publickey_row[782] = `CIPHERTEXT_WIDTH'd15818711;
publickey_row[783] = `CIPHERTEXT_WIDTH'd1955972;
publickey_row[784] = `CIPHERTEXT_WIDTH'd9876255;
publickey_row[785] = `CIPHERTEXT_WIDTH'd6630618;
publickey_row[786] = `CIPHERTEXT_WIDTH'd2578809;
publickey_row[787] = `CIPHERTEXT_WIDTH'd8348399;
publickey_row[788] = `CIPHERTEXT_WIDTH'd5414300;
publickey_row[789] = `CIPHERTEXT_WIDTH'd15833319;
publickey_row[790] = `CIPHERTEXT_WIDTH'd11636034;
publickey_row[791] = `CIPHERTEXT_WIDTH'd1782550;
publickey_row[792] = `CIPHERTEXT_WIDTH'd3091905;
publickey_row[793] = `CIPHERTEXT_WIDTH'd12846082;
publickey_row[794] = `CIPHERTEXT_WIDTH'd15174215;
publickey_row[795] = `CIPHERTEXT_WIDTH'd5495809;
publickey_row[796] = `CIPHERTEXT_WIDTH'd2925177;
publickey_row[797] = `CIPHERTEXT_WIDTH'd822628;
publickey_row[798] = `CIPHERTEXT_WIDTH'd3009926;
publickey_row[799] = `CIPHERTEXT_WIDTH'd15572469;
publickey_row[800] = `CIPHERTEXT_WIDTH'd998638;
publickey_row[801] = `CIPHERTEXT_WIDTH'd8007309;
publickey_row[802] = `CIPHERTEXT_WIDTH'd3158604;
publickey_row[803] = `CIPHERTEXT_WIDTH'd16544062;
publickey_row[804] = `CIPHERTEXT_WIDTH'd1933892;
publickey_row[805] = `CIPHERTEXT_WIDTH'd9837991;
publickey_row[806] = `CIPHERTEXT_WIDTH'd8871850;
publickey_row[807] = `CIPHERTEXT_WIDTH'd16302837;
publickey_row[808] = `CIPHERTEXT_WIDTH'd14373031;
publickey_row[809] = `CIPHERTEXT_WIDTH'd4607250;
publickey_row[810] = `CIPHERTEXT_WIDTH'd14685985;
publickey_row[811] = `CIPHERTEXT_WIDTH'd1693330;
publickey_row[812] = `CIPHERTEXT_WIDTH'd10161618;
publickey_row[813] = `CIPHERTEXT_WIDTH'd11240929;
publickey_row[814] = `CIPHERTEXT_WIDTH'd1138895;
publickey_row[815] = `CIPHERTEXT_WIDTH'd1396358;
publickey_row[816] = `CIPHERTEXT_WIDTH'd11756055;
publickey_row[817] = `CIPHERTEXT_WIDTH'd6855958;
publickey_row[818] = `CIPHERTEXT_WIDTH'd3720635;
publickey_row[819] = `CIPHERTEXT_WIDTH'd13631703;
publickey_row[820] = `CIPHERTEXT_WIDTH'd4441374;
publickey_row[821] = `CIPHERTEXT_WIDTH'd12862530;
publickey_row[822] = `CIPHERTEXT_WIDTH'd7428043;
publickey_row[823] = `CIPHERTEXT_WIDTH'd16639893;
publickey_row[824] = `CIPHERTEXT_WIDTH'd2585917;
publickey_row[825] = `CIPHERTEXT_WIDTH'd13256984;
publickey_row[826] = `CIPHERTEXT_WIDTH'd11071758;
publickey_row[827] = `CIPHERTEXT_WIDTH'd14072672;
publickey_row[828] = `CIPHERTEXT_WIDTH'd4370360;
publickey_row[829] = `CIPHERTEXT_WIDTH'd3662180;
publickey_row[830] = `CIPHERTEXT_WIDTH'd4668010;
publickey_row[831] = `CIPHERTEXT_WIDTH'd7060952;
publickey_row[832] = `CIPHERTEXT_WIDTH'd1623076;
publickey_row[833] = `CIPHERTEXT_WIDTH'd12681782;
publickey_row[834] = `CIPHERTEXT_WIDTH'd3292835;
publickey_row[835] = `CIPHERTEXT_WIDTH'd6760233;
publickey_row[836] = `CIPHERTEXT_WIDTH'd8766396;
publickey_row[837] = `CIPHERTEXT_WIDTH'd16084606;
publickey_row[838] = `CIPHERTEXT_WIDTH'd12809089;
publickey_row[839] = `CIPHERTEXT_WIDTH'd14045839;
publickey_row[840] = `CIPHERTEXT_WIDTH'd11621101;
publickey_row[841] = `CIPHERTEXT_WIDTH'd1828566;
publickey_row[842] = `CIPHERTEXT_WIDTH'd3745557;
publickey_row[843] = `CIPHERTEXT_WIDTH'd10012870;
publickey_row[844] = `CIPHERTEXT_WIDTH'd15004478;
publickey_row[845] = `CIPHERTEXT_WIDTH'd12422879;
publickey_row[846] = `CIPHERTEXT_WIDTH'd6228067;
publickey_row[847] = `CIPHERTEXT_WIDTH'd1093065;
publickey_row[848] = `CIPHERTEXT_WIDTH'd7642992;
publickey_row[849] = `CIPHERTEXT_WIDTH'd12690354;
publickey_row[850] = `CIPHERTEXT_WIDTH'd12239433;
publickey_row[851] = `CIPHERTEXT_WIDTH'd16690619;
publickey_row[852] = `CIPHERTEXT_WIDTH'd9443891;
publickey_row[853] = `CIPHERTEXT_WIDTH'd11138280;
publickey_row[854] = `CIPHERTEXT_WIDTH'd13680100;
publickey_row[855] = `CIPHERTEXT_WIDTH'd281298;
publickey_row[856] = `CIPHERTEXT_WIDTH'd13579994;
publickey_row[857] = `CIPHERTEXT_WIDTH'd13217636;
publickey_row[858] = `CIPHERTEXT_WIDTH'd14232982;
publickey_row[859] = `CIPHERTEXT_WIDTH'd3534487;
publickey_row[860] = `CIPHERTEXT_WIDTH'd14840559;
publickey_row[861] = `CIPHERTEXT_WIDTH'd2845177;
publickey_row[862] = `CIPHERTEXT_WIDTH'd16744433;
publickey_row[863] = `CIPHERTEXT_WIDTH'd11687451;
publickey_row[864] = `CIPHERTEXT_WIDTH'd14504160;
publickey_row[865] = `CIPHERTEXT_WIDTH'd11396987;
publickey_row[866] = `CIPHERTEXT_WIDTH'd783347;
publickey_row[867] = `CIPHERTEXT_WIDTH'd8480652;
publickey_row[868] = `CIPHERTEXT_WIDTH'd14392152;
publickey_row[869] = `CIPHERTEXT_WIDTH'd1257463;
publickey_row[870] = `CIPHERTEXT_WIDTH'd12190539;
publickey_row[871] = `CIPHERTEXT_WIDTH'd1266069;
publickey_row[872] = `CIPHERTEXT_WIDTH'd3057838;
publickey_row[873] = `CIPHERTEXT_WIDTH'd14527402;
publickey_row[874] = `CIPHERTEXT_WIDTH'd1403523;
publickey_row[875] = `CIPHERTEXT_WIDTH'd904584;
publickey_row[876] = `CIPHERTEXT_WIDTH'd2946365;
publickey_row[877] = `CIPHERTEXT_WIDTH'd12451839;
publickey_row[878] = `CIPHERTEXT_WIDTH'd11408264;
publickey_row[879] = `CIPHERTEXT_WIDTH'd1089603;
publickey_row[880] = `CIPHERTEXT_WIDTH'd3160314;
publickey_row[881] = `CIPHERTEXT_WIDTH'd11533152;
publickey_row[882] = `CIPHERTEXT_WIDTH'd10503822;
publickey_row[883] = `CIPHERTEXT_WIDTH'd9055551;
publickey_row[884] = `CIPHERTEXT_WIDTH'd13065781;
publickey_row[885] = `CIPHERTEXT_WIDTH'd10239536;
publickey_row[886] = `CIPHERTEXT_WIDTH'd15767827;
publickey_row[887] = `CIPHERTEXT_WIDTH'd11449549;
publickey_row[888] = `CIPHERTEXT_WIDTH'd9434696;
publickey_row[889] = `CIPHERTEXT_WIDTH'd15181408;
publickey_row[890] = `CIPHERTEXT_WIDTH'd3124137;
publickey_row[891] = `CIPHERTEXT_WIDTH'd8482681;
publickey_row[892] = `CIPHERTEXT_WIDTH'd11543992;
publickey_row[893] = `CIPHERTEXT_WIDTH'd8508119;
publickey_row[894] = `CIPHERTEXT_WIDTH'd11183332;
publickey_row[895] = `CIPHERTEXT_WIDTH'd13468276;
publickey_row[896] = `CIPHERTEXT_WIDTH'd14233600;
publickey_row[897] = `CIPHERTEXT_WIDTH'd1743722;
publickey_row[898] = `CIPHERTEXT_WIDTH'd14385388;
publickey_row[899] = `CIPHERTEXT_WIDTH'd9042170;
publickey_row[900] = `CIPHERTEXT_WIDTH'd10015302;
publickey_row[901] = `CIPHERTEXT_WIDTH'd15914802;
publickey_row[902] = `CIPHERTEXT_WIDTH'd6850584;
publickey_row[903] = `CIPHERTEXT_WIDTH'd986807;
publickey_row[904] = `CIPHERTEXT_WIDTH'd14790346;
publickey_row[905] = `CIPHERTEXT_WIDTH'd2854876;
publickey_row[906] = `CIPHERTEXT_WIDTH'd3288726;
publickey_row[907] = `CIPHERTEXT_WIDTH'd8257253;
publickey_row[908] = `CIPHERTEXT_WIDTH'd9774517;
publickey_row[909] = `CIPHERTEXT_WIDTH'd11878892;
publickey_row[910] = `CIPHERTEXT_WIDTH'd5656076;
publickey_row[911] = `CIPHERTEXT_WIDTH'd1386866;
publickey_row[912] = `CIPHERTEXT_WIDTH'd8484433;
publickey_row[913] = `CIPHERTEXT_WIDTH'd16336234;
publickey_row[914] = `CIPHERTEXT_WIDTH'd10185253;
publickey_row[915] = `CIPHERTEXT_WIDTH'd39260;
publickey_row[916] = `CIPHERTEXT_WIDTH'd3984365;
publickey_row[917] = `CIPHERTEXT_WIDTH'd15439710;
publickey_row[918] = `CIPHERTEXT_WIDTH'd6842915;
publickey_row[919] = `CIPHERTEXT_WIDTH'd12154620;
publickey_row[920] = `CIPHERTEXT_WIDTH'd10486119;
publickey_row[921] = `CIPHERTEXT_WIDTH'd4846804;
publickey_row[922] = `CIPHERTEXT_WIDTH'd14456856;
publickey_row[923] = `CIPHERTEXT_WIDTH'd11409518;
publickey_row[924] = `CIPHERTEXT_WIDTH'd11735954;
publickey_row[925] = `CIPHERTEXT_WIDTH'd12990449;
publickey_row[926] = `CIPHERTEXT_WIDTH'd10567683;
publickey_row[927] = `CIPHERTEXT_WIDTH'd4388728;
publickey_row[928] = `CIPHERTEXT_WIDTH'd10070134;
publickey_row[929] = `CIPHERTEXT_WIDTH'd4622367;
publickey_row[930] = `CIPHERTEXT_WIDTH'd7765653;
publickey_row[931] = `CIPHERTEXT_WIDTH'd7700232;
publickey_row[932] = `CIPHERTEXT_WIDTH'd1608650;
publickey_row[933] = `CIPHERTEXT_WIDTH'd12890024;
publickey_row[934] = `CIPHERTEXT_WIDTH'd1758100;
publickey_row[935] = `CIPHERTEXT_WIDTH'd10139495;
publickey_row[936] = `CIPHERTEXT_WIDTH'd11922465;
publickey_row[937] = `CIPHERTEXT_WIDTH'd9002075;
publickey_row[938] = `CIPHERTEXT_WIDTH'd5215926;
publickey_row[939] = `CIPHERTEXT_WIDTH'd13646754;
publickey_row[940] = `CIPHERTEXT_WIDTH'd2135823;
publickey_row[941] = `CIPHERTEXT_WIDTH'd748423;
publickey_row[942] = `CIPHERTEXT_WIDTH'd5582709;
publickey_row[943] = `CIPHERTEXT_WIDTH'd11250617;
publickey_row[944] = `CIPHERTEXT_WIDTH'd8936549;
publickey_row[945] = `CIPHERTEXT_WIDTH'd5638265;
publickey_row[946] = `CIPHERTEXT_WIDTH'd14241247;
publickey_row[947] = `CIPHERTEXT_WIDTH'd13847396;
publickey_row[948] = `CIPHERTEXT_WIDTH'd13306367;
publickey_row[949] = `CIPHERTEXT_WIDTH'd5641986;
publickey_row[950] = `CIPHERTEXT_WIDTH'd7094205;
publickey_row[951] = `CIPHERTEXT_WIDTH'd11172370;
publickey_row[952] = `CIPHERTEXT_WIDTH'd16404225;
publickey_row[953] = `CIPHERTEXT_WIDTH'd12211381;
publickey_row[954] = `CIPHERTEXT_WIDTH'd1561212;
publickey_row[955] = `CIPHERTEXT_WIDTH'd11140844;
publickey_row[956] = `CIPHERTEXT_WIDTH'd12613288;
publickey_row[957] = `CIPHERTEXT_WIDTH'd4412725;
publickey_row[958] = `CIPHERTEXT_WIDTH'd4570231;
publickey_row[959] = `CIPHERTEXT_WIDTH'd8574941;
publickey_row[960] = `CIPHERTEXT_WIDTH'd7597586;
publickey_row[961] = `CIPHERTEXT_WIDTH'd2451505;
publickey_row[962] = `CIPHERTEXT_WIDTH'd2034390;
publickey_row[963] = `CIPHERTEXT_WIDTH'd16273049;
publickey_row[964] = `CIPHERTEXT_WIDTH'd10333928;
publickey_row[965] = `CIPHERTEXT_WIDTH'd15749407;
publickey_row[966] = `CIPHERTEXT_WIDTH'd10916802;
publickey_row[967] = `CIPHERTEXT_WIDTH'd5145601;
publickey_row[968] = `CIPHERTEXT_WIDTH'd2481552;
publickey_row[969] = `CIPHERTEXT_WIDTH'd8679474;
publickey_row[970] = `CIPHERTEXT_WIDTH'd9550863;
publickey_row[971] = `CIPHERTEXT_WIDTH'd1595961;
publickey_row[972] = `CIPHERTEXT_WIDTH'd2716585;
publickey_row[973] = `CIPHERTEXT_WIDTH'd13476321;
publickey_row[974] = `CIPHERTEXT_WIDTH'd10824225;
publickey_row[975] = `CIPHERTEXT_WIDTH'd3779787;
publickey_row[976] = `CIPHERTEXT_WIDTH'd9788590;
publickey_row[977] = `CIPHERTEXT_WIDTH'd5985231;
publickey_row[978] = `CIPHERTEXT_WIDTH'd2027920;
publickey_row[979] = `CIPHERTEXT_WIDTH'd5479136;
publickey_row[980] = `CIPHERTEXT_WIDTH'd13149374;
publickey_row[981] = `CIPHERTEXT_WIDTH'd10196834;
publickey_row[982] = `CIPHERTEXT_WIDTH'd27773;
publickey_row[983] = `CIPHERTEXT_WIDTH'd7166638;
publickey_row[984] = `CIPHERTEXT_WIDTH'd16457334;
publickey_row[985] = `CIPHERTEXT_WIDTH'd10137377;
publickey_row[986] = `CIPHERTEXT_WIDTH'd13730625;
publickey_row[987] = `CIPHERTEXT_WIDTH'd3043191;
publickey_row[988] = `CIPHERTEXT_WIDTH'd7724325;
publickey_row[989] = `CIPHERTEXT_WIDTH'd14166363;
publickey_row[990] = `CIPHERTEXT_WIDTH'd10802516;
publickey_row[991] = `CIPHERTEXT_WIDTH'd1990443;
publickey_row[992] = `CIPHERTEXT_WIDTH'd999332;
publickey_row[993] = `CIPHERTEXT_WIDTH'd12240946;
publickey_row[994] = `CIPHERTEXT_WIDTH'd7579996;
publickey_row[995] = `CIPHERTEXT_WIDTH'd7474257;
publickey_row[996] = `CIPHERTEXT_WIDTH'd2456188;
publickey_row[997] = `CIPHERTEXT_WIDTH'd7489889;
publickey_row[998] = `CIPHERTEXT_WIDTH'd15102249;
publickey_row[999] = `CIPHERTEXT_WIDTH'd597436;
publickey_row[1000] = `CIPHERTEXT_WIDTH'd15747622;
publickey_row[1001] = `CIPHERTEXT_WIDTH'd11436739;
publickey_row[1002] = `CIPHERTEXT_WIDTH'd6908164;
publickey_row[1003] = `CIPHERTEXT_WIDTH'd3584396;
publickey_row[1004] = `CIPHERTEXT_WIDTH'd15755328;
publickey_row[1005] = `CIPHERTEXT_WIDTH'd10738885;
publickey_row[1006] = `CIPHERTEXT_WIDTH'd10686935;
publickey_row[1007] = `CIPHERTEXT_WIDTH'd9248129;
publickey_row[1008] = `CIPHERTEXT_WIDTH'd2267483;
publickey_row[1009] = `CIPHERTEXT_WIDTH'd224710;
publickey_row[1010] = `CIPHERTEXT_WIDTH'd5430184;
publickey_row[1011] = `CIPHERTEXT_WIDTH'd3291045;
publickey_row[1012] = `CIPHERTEXT_WIDTH'd6580269;
publickey_row[1013] = `CIPHERTEXT_WIDTH'd16581558;
publickey_row[1014] = `CIPHERTEXT_WIDTH'd11069453;
publickey_row[1015] = `CIPHERTEXT_WIDTH'd5296518;
publickey_row[1016] = `CIPHERTEXT_WIDTH'd9825727;
publickey_row[1017] = `CIPHERTEXT_WIDTH'd9497745;
publickey_row[1018] = `CIPHERTEXT_WIDTH'd1615396;
publickey_row[1019] = `CIPHERTEXT_WIDTH'd9146480;
publickey_row[1020] = `CIPHERTEXT_WIDTH'd566885;
publickey_row[1021] = `CIPHERTEXT_WIDTH'd8265970;
publickey_row[1022] = `CIPHERTEXT_WIDTH'd14293051;
publickey_row[1023] = `CIPHERTEXT_WIDTH'd14995949;
publickey_row[1024] = `CIPHERTEXT_WIDTH'd16409631;
publickey_row[1025] = `CIPHERTEXT_WIDTH'd16202846;
publickey_row[1026] = `CIPHERTEXT_WIDTH'd11417742;
publickey_row[1027] = `CIPHERTEXT_WIDTH'd5692406;
publickey_row[1028] = `CIPHERTEXT_WIDTH'd9267784;
publickey_row[1029] = `CIPHERTEXT_WIDTH'd14776342;
publickey_row[1030] = `CIPHERTEXT_WIDTH'd6214245;
publickey_row[1031] = `CIPHERTEXT_WIDTH'd7498942;
publickey_row[1032] = `CIPHERTEXT_WIDTH'd355315;
publickey_row[1033] = `CIPHERTEXT_WIDTH'd773942;
publickey_row[1034] = `CIPHERTEXT_WIDTH'd9534680;
publickey_row[1035] = `CIPHERTEXT_WIDTH'd16733985;
publickey_row[1036] = `CIPHERTEXT_WIDTH'd7647893;
publickey_row[1037] = `CIPHERTEXT_WIDTH'd9958645;
publickey_row[1038] = `CIPHERTEXT_WIDTH'd5258266;
publickey_row[1039] = `CIPHERTEXT_WIDTH'd9515338;
publickey_row[1040] = `CIPHERTEXT_WIDTH'd13168102;
publickey_row[1041] = `CIPHERTEXT_WIDTH'd1619990;
publickey_row[1042] = `CIPHERTEXT_WIDTH'd13367556;
publickey_row[1043] = `CIPHERTEXT_WIDTH'd8204815;
publickey_row[1044] = `CIPHERTEXT_WIDTH'd9506915;
publickey_row[1045] = `CIPHERTEXT_WIDTH'd2445154;
publickey_row[1046] = `CIPHERTEXT_WIDTH'd4869912;
publickey_row[1047] = `CIPHERTEXT_WIDTH'd2311315;
publickey_row[1048] = `CIPHERTEXT_WIDTH'd10252796;
publickey_row[1049] = `CIPHERTEXT_WIDTH'd3232974;
publickey_row[1050] = `CIPHERTEXT_WIDTH'd10140555;
publickey_row[1051] = `CIPHERTEXT_WIDTH'd4358310;
publickey_row[1052] = `CIPHERTEXT_WIDTH'd806554;
publickey_row[1053] = `CIPHERTEXT_WIDTH'd4301044;
publickey_row[1054] = `CIPHERTEXT_WIDTH'd4449760;
publickey_row[1055] = `CIPHERTEXT_WIDTH'd11387505;
publickey_row[1056] = `CIPHERTEXT_WIDTH'd16408465;
publickey_row[1057] = `CIPHERTEXT_WIDTH'd5277676;
publickey_row[1058] = `CIPHERTEXT_WIDTH'd13445891;
publickey_row[1059] = `CIPHERTEXT_WIDTH'd15643121;
publickey_row[1060] = `CIPHERTEXT_WIDTH'd10909933;
publickey_row[1061] = `CIPHERTEXT_WIDTH'd7291347;
publickey_row[1062] = `CIPHERTEXT_WIDTH'd10003825;
publickey_row[1063] = `CIPHERTEXT_WIDTH'd4953370;
publickey_row[1064] = `CIPHERTEXT_WIDTH'd5002190;
publickey_row[1065] = `CIPHERTEXT_WIDTH'd2691540;
publickey_row[1066] = `CIPHERTEXT_WIDTH'd971649;
publickey_row[1067] = `CIPHERTEXT_WIDTH'd1471272;
publickey_row[1068] = `CIPHERTEXT_WIDTH'd351721;
publickey_row[1069] = `CIPHERTEXT_WIDTH'd7914711;
publickey_row[1070] = `CIPHERTEXT_WIDTH'd13560157;
publickey_row[1071] = `CIPHERTEXT_WIDTH'd548114;
publickey_row[1072] = `CIPHERTEXT_WIDTH'd11723488;
publickey_row[1073] = `CIPHERTEXT_WIDTH'd4068750;
publickey_row[1074] = `CIPHERTEXT_WIDTH'd16730070;
publickey_row[1075] = `CIPHERTEXT_WIDTH'd4910284;
publickey_row[1076] = `CIPHERTEXT_WIDTH'd2421536;
publickey_row[1077] = `CIPHERTEXT_WIDTH'd3507826;
publickey_row[1078] = `CIPHERTEXT_WIDTH'd13880968;
publickey_row[1079] = `CIPHERTEXT_WIDTH'd6050292;
publickey_row[1080] = `CIPHERTEXT_WIDTH'd10433200;
publickey_row[1081] = `CIPHERTEXT_WIDTH'd1107774;
publickey_row[1082] = `CIPHERTEXT_WIDTH'd15448797;
publickey_row[1083] = `CIPHERTEXT_WIDTH'd13067381;
publickey_row[1084] = `CIPHERTEXT_WIDTH'd2669404;
publickey_row[1085] = `CIPHERTEXT_WIDTH'd13658022;
publickey_row[1086] = `CIPHERTEXT_WIDTH'd15020874;
publickey_row[1087] = `CIPHERTEXT_WIDTH'd2566355;
publickey_row[1088] = `CIPHERTEXT_WIDTH'd9518663;
publickey_row[1089] = `CIPHERTEXT_WIDTH'd12376427;
publickey_row[1090] = `CIPHERTEXT_WIDTH'd1706882;
publickey_row[1091] = `CIPHERTEXT_WIDTH'd2235313;
publickey_row[1092] = `CIPHERTEXT_WIDTH'd7439247;
publickey_row[1093] = `CIPHERTEXT_WIDTH'd13867643;
publickey_row[1094] = `CIPHERTEXT_WIDTH'd12687371;
publickey_row[1095] = `CIPHERTEXT_WIDTH'd10439137;
publickey_row[1096] = `CIPHERTEXT_WIDTH'd9110189;
publickey_row[1097] = `CIPHERTEXT_WIDTH'd4398087;
publickey_row[1098] = `CIPHERTEXT_WIDTH'd12465809;
publickey_row[1099] = `CIPHERTEXT_WIDTH'd5187051;
publickey_row[1100] = `CIPHERTEXT_WIDTH'd13878600;
publickey_row[1101] = `CIPHERTEXT_WIDTH'd7646833;
publickey_row[1102] = `CIPHERTEXT_WIDTH'd4533946;
publickey_row[1103] = `CIPHERTEXT_WIDTH'd7411241;
publickey_row[1104] = `CIPHERTEXT_WIDTH'd11138564;
publickey_row[1105] = `CIPHERTEXT_WIDTH'd3802883;
publickey_row[1106] = `CIPHERTEXT_WIDTH'd8900862;
publickey_row[1107] = `CIPHERTEXT_WIDTH'd11871203;
publickey_row[1108] = `CIPHERTEXT_WIDTH'd11948455;
publickey_row[1109] = `CIPHERTEXT_WIDTH'd8612993;
publickey_row[1110] = `CIPHERTEXT_WIDTH'd8493146;
publickey_row[1111] = `CIPHERTEXT_WIDTH'd2561286;
publickey_row[1112] = `CIPHERTEXT_WIDTH'd14720447;
publickey_row[1113] = `CIPHERTEXT_WIDTH'd7164988;
publickey_row[1114] = `CIPHERTEXT_WIDTH'd13085318;
publickey_row[1115] = `CIPHERTEXT_WIDTH'd12983057;
publickey_row[1116] = `CIPHERTEXT_WIDTH'd8434006;
publickey_row[1117] = `CIPHERTEXT_WIDTH'd2827564;
publickey_row[1118] = `CIPHERTEXT_WIDTH'd1519161;
publickey_row[1119] = `CIPHERTEXT_WIDTH'd9256110;
publickey_row[1120] = `CIPHERTEXT_WIDTH'd10299083;
publickey_row[1121] = `CIPHERTEXT_WIDTH'd4266559;
publickey_row[1122] = `CIPHERTEXT_WIDTH'd11594276;
publickey_row[1123] = `CIPHERTEXT_WIDTH'd2778581;
publickey_row[1124] = `CIPHERTEXT_WIDTH'd16034890;
publickey_row[1125] = `CIPHERTEXT_WIDTH'd4386759;
publickey_row[1126] = `CIPHERTEXT_WIDTH'd10689904;
publickey_row[1127] = `CIPHERTEXT_WIDTH'd16641859;
publickey_row[1128] = `CIPHERTEXT_WIDTH'd555680;
publickey_row[1129] = `CIPHERTEXT_WIDTH'd8809735;
publickey_row[1130] = `CIPHERTEXT_WIDTH'd3102897;
publickey_row[1131] = `CIPHERTEXT_WIDTH'd4963070;
publickey_row[1132] = `CIPHERTEXT_WIDTH'd2463044;
publickey_row[1133] = `CIPHERTEXT_WIDTH'd11367145;
publickey_row[1134] = `CIPHERTEXT_WIDTH'd2836745;
publickey_row[1135] = `CIPHERTEXT_WIDTH'd2441584;
publickey_row[1136] = `CIPHERTEXT_WIDTH'd11222238;
publickey_row[1137] = `CIPHERTEXT_WIDTH'd15199622;
publickey_row[1138] = `CIPHERTEXT_WIDTH'd15805868;
publickey_row[1139] = `CIPHERTEXT_WIDTH'd13524239;
publickey_row[1140] = `CIPHERTEXT_WIDTH'd16454105;
publickey_row[1141] = `CIPHERTEXT_WIDTH'd7462625;
publickey_row[1142] = `CIPHERTEXT_WIDTH'd8086865;
publickey_row[1143] = `CIPHERTEXT_WIDTH'd1622608;
publickey_row[1144] = `CIPHERTEXT_WIDTH'd8194029;
publickey_row[1145] = `CIPHERTEXT_WIDTH'd16174397;
publickey_row[1146] = `CIPHERTEXT_WIDTH'd15315450;
publickey_row[1147] = `CIPHERTEXT_WIDTH'd16649737;
publickey_row[1148] = `CIPHERTEXT_WIDTH'd1864708;
publickey_row[1149] = `CIPHERTEXT_WIDTH'd679540;
publickey_row[1150] = `CIPHERTEXT_WIDTH'd786590;
publickey_row[1151] = `CIPHERTEXT_WIDTH'd16395713;
publickey_row[1152] = `CIPHERTEXT_WIDTH'd13174097;
publickey_row[1153] = `CIPHERTEXT_WIDTH'd2665134;
publickey_row[1154] = `CIPHERTEXT_WIDTH'd7959756;
publickey_row[1155] = `CIPHERTEXT_WIDTH'd10783491;
publickey_row[1156] = `CIPHERTEXT_WIDTH'd9645841;
publickey_row[1157] = `CIPHERTEXT_WIDTH'd14320893;
publickey_row[1158] = `CIPHERTEXT_WIDTH'd3360309;
publickey_row[1159] = `CIPHERTEXT_WIDTH'd5779718;
publickey_row[1160] = `CIPHERTEXT_WIDTH'd16504968;
publickey_row[1161] = `CIPHERTEXT_WIDTH'd10319051;
publickey_row[1162] = `CIPHERTEXT_WIDTH'd15558634;
publickey_row[1163] = `CIPHERTEXT_WIDTH'd5620205;
publickey_row[1164] = `CIPHERTEXT_WIDTH'd718508;
publickey_row[1165] = `CIPHERTEXT_WIDTH'd3976404;
publickey_row[1166] = `CIPHERTEXT_WIDTH'd10517751;
publickey_row[1167] = `CIPHERTEXT_WIDTH'd11487709;
publickey_row[1168] = `CIPHERTEXT_WIDTH'd11709404;
publickey_row[1169] = `CIPHERTEXT_WIDTH'd1635809;
publickey_row[1170] = `CIPHERTEXT_WIDTH'd3668832;
publickey_row[1171] = `CIPHERTEXT_WIDTH'd7846343;
publickey_row[1172] = `CIPHERTEXT_WIDTH'd16462445;
publickey_row[1173] = `CIPHERTEXT_WIDTH'd13346979;
publickey_row[1174] = `CIPHERTEXT_WIDTH'd11601870;
publickey_row[1175] = `CIPHERTEXT_WIDTH'd16270123;
publickey_row[1176] = `CIPHERTEXT_WIDTH'd1934169;
publickey_row[1177] = `CIPHERTEXT_WIDTH'd4310472;
publickey_row[1178] = `CIPHERTEXT_WIDTH'd4872426;
publickey_row[1179] = `CIPHERTEXT_WIDTH'd9380958;
publickey_row[1180] = `CIPHERTEXT_WIDTH'd450331;
publickey_row[1181] = `CIPHERTEXT_WIDTH'd16359916;
publickey_row[1182] = `CIPHERTEXT_WIDTH'd8090882;
publickey_row[1183] = `CIPHERTEXT_WIDTH'd4732297;
publickey_row[1184] = `CIPHERTEXT_WIDTH'd6067613;
publickey_row[1185] = `CIPHERTEXT_WIDTH'd10181944;
publickey_row[1186] = `CIPHERTEXT_WIDTH'd6000441;
publickey_row[1187] = `CIPHERTEXT_WIDTH'd10800252;
publickey_row[1188] = `CIPHERTEXT_WIDTH'd2606996;
publickey_row[1189] = `CIPHERTEXT_WIDTH'd15022668;
publickey_row[1190] = `CIPHERTEXT_WIDTH'd7960704;
publickey_row[1191] = `CIPHERTEXT_WIDTH'd4816142;
publickey_row[1192] = `CIPHERTEXT_WIDTH'd9349034;
publickey_row[1193] = `CIPHERTEXT_WIDTH'd14179825;
publickey_row[1194] = `CIPHERTEXT_WIDTH'd10291335;
publickey_row[1195] = `CIPHERTEXT_WIDTH'd3236846;
publickey_row[1196] = `CIPHERTEXT_WIDTH'd2550906;
publickey_row[1197] = `CIPHERTEXT_WIDTH'd5218625;
publickey_row[1198] = `CIPHERTEXT_WIDTH'd2046593;
publickey_row[1199] = `CIPHERTEXT_WIDTH'd9499313;
publickey_row[1200] = `CIPHERTEXT_WIDTH'd15694943;
publickey_row[1201] = `CIPHERTEXT_WIDTH'd11215181;
publickey_row[1202] = `CIPHERTEXT_WIDTH'd15648525;
publickey_row[1203] = `CIPHERTEXT_WIDTH'd6269468;
publickey_row[1204] = `CIPHERTEXT_WIDTH'd5802850;
publickey_row[1205] = `CIPHERTEXT_WIDTH'd5687698;
publickey_row[1206] = `CIPHERTEXT_WIDTH'd3417580;
publickey_row[1207] = `CIPHERTEXT_WIDTH'd10151656;
publickey_row[1208] = `CIPHERTEXT_WIDTH'd2183794;
publickey_row[1209] = `CIPHERTEXT_WIDTH'd14340483;
publickey_row[1210] = `CIPHERTEXT_WIDTH'd13110585;
publickey_row[1211] = `CIPHERTEXT_WIDTH'd9274834;
publickey_row[1212] = `CIPHERTEXT_WIDTH'd12734694;
publickey_row[1213] = `CIPHERTEXT_WIDTH'd3805416;
publickey_row[1214] = `CIPHERTEXT_WIDTH'd1423067;
publickey_row[1215] = `CIPHERTEXT_WIDTH'd9271190;
publickey_row[1216] = `CIPHERTEXT_WIDTH'd12536221;
publickey_row[1217] = `CIPHERTEXT_WIDTH'd1904847;
publickey_row[1218] = `CIPHERTEXT_WIDTH'd12713864;
publickey_row[1219] = `CIPHERTEXT_WIDTH'd1309086;
publickey_row[1220] = `CIPHERTEXT_WIDTH'd64634;
publickey_row[1221] = `CIPHERTEXT_WIDTH'd11105279;
publickey_row[1222] = `CIPHERTEXT_WIDTH'd2340609;
publickey_row[1223] = `CIPHERTEXT_WIDTH'd1496307;
publickey_row[1224] = `CIPHERTEXT_WIDTH'd6512379;
publickey_row[1225] = `CIPHERTEXT_WIDTH'd2898588;
publickey_row[1226] = `CIPHERTEXT_WIDTH'd9810387;
publickey_row[1227] = `CIPHERTEXT_WIDTH'd8053046;
publickey_row[1228] = `CIPHERTEXT_WIDTH'd7334212;
publickey_row[1229] = `CIPHERTEXT_WIDTH'd142078;
publickey_row[1230] = `CIPHERTEXT_WIDTH'd7195016;
publickey_row[1231] = `CIPHERTEXT_WIDTH'd4435368;
publickey_row[1232] = `CIPHERTEXT_WIDTH'd10725852;
publickey_row[1233] = `CIPHERTEXT_WIDTH'd9348201;
publickey_row[1234] = `CIPHERTEXT_WIDTH'd13266914;
publickey_row[1235] = `CIPHERTEXT_WIDTH'd5676692;
publickey_row[1236] = `CIPHERTEXT_WIDTH'd3500705;
publickey_row[1237] = `CIPHERTEXT_WIDTH'd3940200;
publickey_row[1238] = `CIPHERTEXT_WIDTH'd11135797;
publickey_row[1239] = `CIPHERTEXT_WIDTH'd10287369;
publickey_row[1240] = `CIPHERTEXT_WIDTH'd5624099;
publickey_row[1241] = `CIPHERTEXT_WIDTH'd15306350;
publickey_row[1242] = `CIPHERTEXT_WIDTH'd15870329;
publickey_row[1243] = `CIPHERTEXT_WIDTH'd14711235;
publickey_row[1244] = `CIPHERTEXT_WIDTH'd1723036;
publickey_row[1245] = `CIPHERTEXT_WIDTH'd7614630;
publickey_row[1246] = `CIPHERTEXT_WIDTH'd1105351;
publickey_row[1247] = `CIPHERTEXT_WIDTH'd9297922;
publickey_row[1248] = `CIPHERTEXT_WIDTH'd2743692;
publickey_row[1249] = `CIPHERTEXT_WIDTH'd3859804;
publickey_row[1250] = `CIPHERTEXT_WIDTH'd2539774;
publickey_row[1251] = `CIPHERTEXT_WIDTH'd9732458;
publickey_row[1252] = `CIPHERTEXT_WIDTH'd13712102;
publickey_row[1253] = `CIPHERTEXT_WIDTH'd12389381;
publickey_row[1254] = `CIPHERTEXT_WIDTH'd12849779;
publickey_row[1255] = `CIPHERTEXT_WIDTH'd9326905;
publickey_row[1256] = `CIPHERTEXT_WIDTH'd15204054;
publickey_row[1257] = `CIPHERTEXT_WIDTH'd6646173;
publickey_row[1258] = `CIPHERTEXT_WIDTH'd5196397;
publickey_row[1259] = `CIPHERTEXT_WIDTH'd15348804;
publickey_row[1260] = `CIPHERTEXT_WIDTH'd2030390;
publickey_row[1261] = `CIPHERTEXT_WIDTH'd16150245;
publickey_row[1262] = `CIPHERTEXT_WIDTH'd7919664;
publickey_row[1263] = `CIPHERTEXT_WIDTH'd10282042;
publickey_row[1264] = `CIPHERTEXT_WIDTH'd16091061;
publickey_row[1265] = `CIPHERTEXT_WIDTH'd16722222;
publickey_row[1266] = `CIPHERTEXT_WIDTH'd14025414;
publickey_row[1267] = `CIPHERTEXT_WIDTH'd8057568;
publickey_row[1268] = `CIPHERTEXT_WIDTH'd1033709;
publickey_row[1269] = `CIPHERTEXT_WIDTH'd1769131;
publickey_row[1270] = `CIPHERTEXT_WIDTH'd4211160;
publickey_row[1271] = `CIPHERTEXT_WIDTH'd11682230;
publickey_row[1272] = `CIPHERTEXT_WIDTH'd14124871;
publickey_row[1273] = `CIPHERTEXT_WIDTH'd16655783;
publickey_row[1274] = `CIPHERTEXT_WIDTH'd328504;
publickey_row[1275] = `CIPHERTEXT_WIDTH'd10749179;
publickey_row[1276] = `CIPHERTEXT_WIDTH'd13078314;
publickey_row[1277] = `CIPHERTEXT_WIDTH'd16052447;
publickey_row[1278] = `CIPHERTEXT_WIDTH'd12316651;
publickey_row[1279] = `CIPHERTEXT_WIDTH'd10498624;
publickey_row[1280] = `CIPHERTEXT_WIDTH'd14654456;
publickey_row[1281] = `CIPHERTEXT_WIDTH'd3144954;
publickey_row[1282] = `CIPHERTEXT_WIDTH'd15397538;
publickey_row[1283] = `CIPHERTEXT_WIDTH'd11191816;
publickey_row[1284] = `CIPHERTEXT_WIDTH'd2981149;
publickey_row[1285] = `CIPHERTEXT_WIDTH'd15082669;
publickey_row[1286] = `CIPHERTEXT_WIDTH'd6553996;
publickey_row[1287] = `CIPHERTEXT_WIDTH'd7037083;
publickey_row[1288] = `CIPHERTEXT_WIDTH'd14971074;
publickey_row[1289] = `CIPHERTEXT_WIDTH'd6375511;
publickey_row[1290] = `CIPHERTEXT_WIDTH'd15503447;
publickey_row[1291] = `CIPHERTEXT_WIDTH'd9712879;
publickey_row[1292] = `CIPHERTEXT_WIDTH'd11883576;
publickey_row[1293] = `CIPHERTEXT_WIDTH'd12422176;
publickey_row[1294] = `CIPHERTEXT_WIDTH'd9411619;
publickey_row[1295] = `CIPHERTEXT_WIDTH'd10565635;
publickey_row[1296] = `CIPHERTEXT_WIDTH'd599955;
publickey_row[1297] = `CIPHERTEXT_WIDTH'd5988849;
publickey_row[1298] = `CIPHERTEXT_WIDTH'd12682897;
publickey_row[1299] = `CIPHERTEXT_WIDTH'd5614574;
publickey_row[1300] = `CIPHERTEXT_WIDTH'd4471231;
publickey_row[1301] = `CIPHERTEXT_WIDTH'd5665164;
publickey_row[1302] = `CIPHERTEXT_WIDTH'd7435037;
publickey_row[1303] = `CIPHERTEXT_WIDTH'd8771186;
publickey_row[1304] = `CIPHERTEXT_WIDTH'd2886269;
publickey_row[1305] = `CIPHERTEXT_WIDTH'd15438997;
publickey_row[1306] = `CIPHERTEXT_WIDTH'd9643114;
publickey_row[1307] = `CIPHERTEXT_WIDTH'd11052713;
publickey_row[1308] = `CIPHERTEXT_WIDTH'd9468640;
publickey_row[1309] = `CIPHERTEXT_WIDTH'd7431248;
publickey_row[1310] = `CIPHERTEXT_WIDTH'd15692825;
publickey_row[1311] = `CIPHERTEXT_WIDTH'd16027780;
publickey_row[1312] = `CIPHERTEXT_WIDTH'd14377538;
publickey_row[1313] = `CIPHERTEXT_WIDTH'd10615130;
publickey_row[1314] = `CIPHERTEXT_WIDTH'd9330908;
publickey_row[1315] = `CIPHERTEXT_WIDTH'd9163995;
publickey_row[1316] = `CIPHERTEXT_WIDTH'd4275829;
publickey_row[1317] = `CIPHERTEXT_WIDTH'd11875970;
publickey_row[1318] = `CIPHERTEXT_WIDTH'd1747986;
publickey_row[1319] = `CIPHERTEXT_WIDTH'd8688343;
publickey_row[1320] = `CIPHERTEXT_WIDTH'd3273100;
publickey_row[1321] = `CIPHERTEXT_WIDTH'd3992033;
publickey_row[1322] = `CIPHERTEXT_WIDTH'd16596048;
publickey_row[1323] = `CIPHERTEXT_WIDTH'd1973863;
publickey_row[1324] = `CIPHERTEXT_WIDTH'd2313139;
publickey_row[1325] = `CIPHERTEXT_WIDTH'd509853;
publickey_row[1326] = `CIPHERTEXT_WIDTH'd6069107;
publickey_row[1327] = `CIPHERTEXT_WIDTH'd14208430;
publickey_row[1328] = `CIPHERTEXT_WIDTH'd8082408;
publickey_row[1329] = `CIPHERTEXT_WIDTH'd6836349;
publickey_row[1330] = `CIPHERTEXT_WIDTH'd4579159;
publickey_row[1331] = `CIPHERTEXT_WIDTH'd5411040;
publickey_row[1332] = `CIPHERTEXT_WIDTH'd4025836;
publickey_row[1333] = `CIPHERTEXT_WIDTH'd5491045;
publickey_row[1334] = `CIPHERTEXT_WIDTH'd12154884;
publickey_row[1335] = `CIPHERTEXT_WIDTH'd6311877;
publickey_row[1336] = `CIPHERTEXT_WIDTH'd8529263;
publickey_row[1337] = `CIPHERTEXT_WIDTH'd8628504;
publickey_row[1338] = `CIPHERTEXT_WIDTH'd10643834;
publickey_row[1339] = `CIPHERTEXT_WIDTH'd2376055;
publickey_row[1340] = `CIPHERTEXT_WIDTH'd6103431;
publickey_row[1341] = `CIPHERTEXT_WIDTH'd7660482;
publickey_row[1342] = `CIPHERTEXT_WIDTH'd13477422;
publickey_row[1343] = `CIPHERTEXT_WIDTH'd6837299;
publickey_row[1344] = `CIPHERTEXT_WIDTH'd14719242;
publickey_row[1345] = `CIPHERTEXT_WIDTH'd4865011;
publickey_row[1346] = `CIPHERTEXT_WIDTH'd482969;
publickey_row[1347] = `CIPHERTEXT_WIDTH'd4215777;
publickey_row[1348] = `CIPHERTEXT_WIDTH'd6822723;
publickey_row[1349] = `CIPHERTEXT_WIDTH'd7880237;
publickey_row[1350] = `CIPHERTEXT_WIDTH'd8141503;
publickey_row[1351] = `CIPHERTEXT_WIDTH'd5798722;
publickey_row[1352] = `CIPHERTEXT_WIDTH'd7000160;
publickey_row[1353] = `CIPHERTEXT_WIDTH'd6035063;
publickey_row[1354] = `CIPHERTEXT_WIDTH'd1449796;
publickey_row[1355] = `CIPHERTEXT_WIDTH'd2400719;
publickey_row[1356] = `CIPHERTEXT_WIDTH'd4510633;
publickey_row[1357] = `CIPHERTEXT_WIDTH'd7609792;
publickey_row[1358] = `CIPHERTEXT_WIDTH'd12947264;
publickey_row[1359] = `CIPHERTEXT_WIDTH'd4574636;
publickey_row[1360] = `CIPHERTEXT_WIDTH'd3104469;
publickey_row[1361] = `CIPHERTEXT_WIDTH'd8760470;
publickey_row[1362] = `CIPHERTEXT_WIDTH'd7459435;
publickey_row[1363] = `CIPHERTEXT_WIDTH'd9996071;
publickey_row[1364] = `CIPHERTEXT_WIDTH'd3269811;
publickey_row[1365] = `CIPHERTEXT_WIDTH'd1696758;
publickey_row[1366] = `CIPHERTEXT_WIDTH'd13108168;
publickey_row[1367] = `CIPHERTEXT_WIDTH'd15571830;
publickey_row[1368] = `CIPHERTEXT_WIDTH'd14059788;
publickey_row[1369] = `CIPHERTEXT_WIDTH'd14420125;
publickey_row[1370] = `CIPHERTEXT_WIDTH'd4559977;
publickey_row[1371] = `CIPHERTEXT_WIDTH'd10876853;
publickey_row[1372] = `CIPHERTEXT_WIDTH'd6032792;
publickey_row[1373] = `CIPHERTEXT_WIDTH'd11934795;
publickey_row[1374] = `CIPHERTEXT_WIDTH'd10133680;
publickey_row[1375] = `CIPHERTEXT_WIDTH'd634595;
publickey_row[1376] = `CIPHERTEXT_WIDTH'd6144800;
publickey_row[1377] = `CIPHERTEXT_WIDTH'd16665199;
publickey_row[1378] = `CIPHERTEXT_WIDTH'd82363;
publickey_row[1379] = `CIPHERTEXT_WIDTH'd2643511;
publickey_row[1380] = `CIPHERTEXT_WIDTH'd56862;
publickey_row[1381] = `CIPHERTEXT_WIDTH'd5113794;
publickey_row[1382] = `CIPHERTEXT_WIDTH'd12404308;
publickey_row[1383] = `CIPHERTEXT_WIDTH'd2977458;
publickey_row[1384] = `CIPHERTEXT_WIDTH'd11635043;
publickey_row[1385] = `CIPHERTEXT_WIDTH'd12823217;
publickey_row[1386] = `CIPHERTEXT_WIDTH'd1520779;
publickey_row[1387] = `CIPHERTEXT_WIDTH'd386479;
publickey_row[1388] = `CIPHERTEXT_WIDTH'd9311362;
publickey_row[1389] = `CIPHERTEXT_WIDTH'd7813205;
publickey_row[1390] = `CIPHERTEXT_WIDTH'd6548674;
publickey_row[1391] = `CIPHERTEXT_WIDTH'd6869505;
publickey_row[1392] = `CIPHERTEXT_WIDTH'd15965397;
publickey_row[1393] = `CIPHERTEXT_WIDTH'd14498635;
publickey_row[1394] = `CIPHERTEXT_WIDTH'd1852058;
publickey_row[1395] = `CIPHERTEXT_WIDTH'd689169;
publickey_row[1396] = `CIPHERTEXT_WIDTH'd8295621;
publickey_row[1397] = `CIPHERTEXT_WIDTH'd11275203;
publickey_row[1398] = `CIPHERTEXT_WIDTH'd1811973;
publickey_row[1399] = `CIPHERTEXT_WIDTH'd9833589;
publickey_row[1400] = `CIPHERTEXT_WIDTH'd8814025;
publickey_row[1401] = `CIPHERTEXT_WIDTH'd15473438;
publickey_row[1402] = `CIPHERTEXT_WIDTH'd14338543;
publickey_row[1403] = `CIPHERTEXT_WIDTH'd9694168;
publickey_row[1404] = `CIPHERTEXT_WIDTH'd7007053;
publickey_row[1405] = `CIPHERTEXT_WIDTH'd12473716;
publickey_row[1406] = `CIPHERTEXT_WIDTH'd6164248;
publickey_row[1407] = `CIPHERTEXT_WIDTH'd4562425;
publickey_row[1408] = `CIPHERTEXT_WIDTH'd221473;
publickey_row[1409] = `CIPHERTEXT_WIDTH'd9052864;
publickey_row[1410] = `CIPHERTEXT_WIDTH'd14642558;
publickey_row[1411] = `CIPHERTEXT_WIDTH'd403661;
publickey_row[1412] = `CIPHERTEXT_WIDTH'd13658770;
publickey_row[1413] = `CIPHERTEXT_WIDTH'd5596148;
publickey_row[1414] = `CIPHERTEXT_WIDTH'd11203503;
publickey_row[1415] = `CIPHERTEXT_WIDTH'd15557949;
publickey_row[1416] = `CIPHERTEXT_WIDTH'd9968135;
publickey_row[1417] = `CIPHERTEXT_WIDTH'd16746549;
publickey_row[1418] = `CIPHERTEXT_WIDTH'd16456201;
publickey_row[1419] = `CIPHERTEXT_WIDTH'd7327620;
publickey_row[1420] = `CIPHERTEXT_WIDTH'd9860048;
publickey_row[1421] = `CIPHERTEXT_WIDTH'd1109408;
publickey_row[1422] = `CIPHERTEXT_WIDTH'd10413517;
publickey_row[1423] = `CIPHERTEXT_WIDTH'd7162143;
publickey_row[1424] = `CIPHERTEXT_WIDTH'd9349937;
publickey_row[1425] = `CIPHERTEXT_WIDTH'd11357676;
publickey_row[1426] = `CIPHERTEXT_WIDTH'd8041198;
publickey_row[1427] = `CIPHERTEXT_WIDTH'd2041483;
publickey_row[1428] = `CIPHERTEXT_WIDTH'd7192591;
publickey_row[1429] = `CIPHERTEXT_WIDTH'd2251498;
publickey_row[1430] = `CIPHERTEXT_WIDTH'd9461411;
publickey_row[1431] = `CIPHERTEXT_WIDTH'd15239084;
publickey_row[1432] = `CIPHERTEXT_WIDTH'd2746801;
publickey_row[1433] = `CIPHERTEXT_WIDTH'd6453324;
publickey_row[1434] = `CIPHERTEXT_WIDTH'd1490333;
publickey_row[1435] = `CIPHERTEXT_WIDTH'd13890989;
publickey_row[1436] = `CIPHERTEXT_WIDTH'd4948709;
publickey_row[1437] = `CIPHERTEXT_WIDTH'd12401296;
publickey_row[1438] = `CIPHERTEXT_WIDTH'd4595821;
publickey_row[1439] = `CIPHERTEXT_WIDTH'd10134428;
publickey_row[1440] = `CIPHERTEXT_WIDTH'd5066173;
publickey_row[1441] = `CIPHERTEXT_WIDTH'd4946804;
publickey_row[1442] = `CIPHERTEXT_WIDTH'd10458029;
publickey_row[1443] = `CIPHERTEXT_WIDTH'd11408994;
publickey_row[1444] = `CIPHERTEXT_WIDTH'd16078615;
publickey_row[1445] = `CIPHERTEXT_WIDTH'd6001884;
publickey_row[1446] = `CIPHERTEXT_WIDTH'd13356366;
publickey_row[1447] = `CIPHERTEXT_WIDTH'd13206206;
publickey_row[1448] = `CIPHERTEXT_WIDTH'd10946836;
publickey_row[1449] = `CIPHERTEXT_WIDTH'd4626149;
publickey_row[1450] = `CIPHERTEXT_WIDTH'd16622612;
publickey_row[1451] = `CIPHERTEXT_WIDTH'd2221500;
publickey_row[1452] = `CIPHERTEXT_WIDTH'd6330980;
publickey_row[1453] = `CIPHERTEXT_WIDTH'd7865678;
publickey_row[1454] = `CIPHERTEXT_WIDTH'd15451781;
publickey_row[1455] = `CIPHERTEXT_WIDTH'd4361013;
publickey_row[1456] = `CIPHERTEXT_WIDTH'd2768988;
publickey_row[1457] = `CIPHERTEXT_WIDTH'd11560994;
publickey_row[1458] = `CIPHERTEXT_WIDTH'd9133257;
publickey_row[1459] = `CIPHERTEXT_WIDTH'd9663501;
publickey_row[1460] = `CIPHERTEXT_WIDTH'd6544740;
publickey_row[1461] = `CIPHERTEXT_WIDTH'd1617885;
publickey_row[1462] = `CIPHERTEXT_WIDTH'd8421033;
publickey_row[1463] = `CIPHERTEXT_WIDTH'd10552933;
publickey_row[1464] = `CIPHERTEXT_WIDTH'd14165919;
publickey_row[1465] = `CIPHERTEXT_WIDTH'd6174714;
publickey_row[1466] = `CIPHERTEXT_WIDTH'd5872272;
publickey_row[1467] = `CIPHERTEXT_WIDTH'd9632570;
publickey_row[1468] = `CIPHERTEXT_WIDTH'd10085399;
publickey_row[1469] = `CIPHERTEXT_WIDTH'd12325580;
publickey_row[1470] = `CIPHERTEXT_WIDTH'd13597975;
publickey_row[1471] = `CIPHERTEXT_WIDTH'd816081;
publickey_row[1472] = `CIPHERTEXT_WIDTH'd12341159;
publickey_row[1473] = `CIPHERTEXT_WIDTH'd13106166;
publickey_row[1474] = `CIPHERTEXT_WIDTH'd6290735;
publickey_row[1475] = `CIPHERTEXT_WIDTH'd12678488;
publickey_row[1476] = `CIPHERTEXT_WIDTH'd9361447;
publickey_row[1477] = `CIPHERTEXT_WIDTH'd12588968;
publickey_row[1478] = `CIPHERTEXT_WIDTH'd9162748;
publickey_row[1479] = `CIPHERTEXT_WIDTH'd1303438;
publickey_row[1480] = `CIPHERTEXT_WIDTH'd645787;
publickey_row[1481] = `CIPHERTEXT_WIDTH'd9511710;
publickey_row[1482] = `CIPHERTEXT_WIDTH'd6130947;
publickey_row[1483] = `CIPHERTEXT_WIDTH'd14379211;
publickey_row[1484] = `CIPHERTEXT_WIDTH'd1448935;
publickey_row[1485] = `CIPHERTEXT_WIDTH'd3822928;
publickey_row[1486] = `CIPHERTEXT_WIDTH'd16399949;
publickey_row[1487] = `CIPHERTEXT_WIDTH'd11702689;
publickey_row[1488] = `CIPHERTEXT_WIDTH'd16576047;
publickey_row[1489] = `CIPHERTEXT_WIDTH'd8422097;
publickey_row[1490] = `CIPHERTEXT_WIDTH'd8366508;
publickey_row[1491] = `CIPHERTEXT_WIDTH'd5030209;
publickey_row[1492] = `CIPHERTEXT_WIDTH'd14752735;
publickey_row[1493] = `CIPHERTEXT_WIDTH'd16425441;
publickey_row[1494] = `CIPHERTEXT_WIDTH'd7510681;
publickey_row[1495] = `CIPHERTEXT_WIDTH'd3110454;
publickey_row[1496] = `CIPHERTEXT_WIDTH'd11949572;
publickey_row[1497] = `CIPHERTEXT_WIDTH'd4839618;
publickey_row[1498] = `CIPHERTEXT_WIDTH'd10740682;
publickey_row[1499] = `CIPHERTEXT_WIDTH'd9718618;
publickey_row[1500] = `CIPHERTEXT_WIDTH'd2139950;
publickey_row[1501] = `CIPHERTEXT_WIDTH'd11805824;
publickey_row[1502] = `CIPHERTEXT_WIDTH'd15004773;
publickey_row[1503] = `CIPHERTEXT_WIDTH'd14395575;
publickey_row[1504] = `CIPHERTEXT_WIDTH'd13727929;
publickey_row[1505] = `CIPHERTEXT_WIDTH'd14843127;
publickey_row[1506] = `CIPHERTEXT_WIDTH'd9343867;
publickey_row[1507] = `CIPHERTEXT_WIDTH'd1301411;
publickey_row[1508] = `CIPHERTEXT_WIDTH'd3012373;
publickey_row[1509] = `CIPHERTEXT_WIDTH'd11959599;
publickey_row[1510] = `CIPHERTEXT_WIDTH'd5067737;
publickey_row[1511] = `CIPHERTEXT_WIDTH'd355149;
publickey_row[1512] = `CIPHERTEXT_WIDTH'd1880297;
publickey_row[1513] = `CIPHERTEXT_WIDTH'd1991323;
publickey_row[1514] = `CIPHERTEXT_WIDTH'd7013634;
publickey_row[1515] = `CIPHERTEXT_WIDTH'd16602193;
publickey_row[1516] = `CIPHERTEXT_WIDTH'd14832517;
publickey_row[1517] = `CIPHERTEXT_WIDTH'd12194781;
publickey_row[1518] = `CIPHERTEXT_WIDTH'd10479511;
publickey_row[1519] = `CIPHERTEXT_WIDTH'd3471290;
publickey_row[1520] = `CIPHERTEXT_WIDTH'd6939253;
publickey_row[1521] = `CIPHERTEXT_WIDTH'd10192381;
publickey_row[1522] = `CIPHERTEXT_WIDTH'd4011981;
publickey_row[1523] = `CIPHERTEXT_WIDTH'd8353218;
publickey_row[1524] = `CIPHERTEXT_WIDTH'd14520584;
publickey_row[1525] = `CIPHERTEXT_WIDTH'd1208962;
publickey_row[1526] = `CIPHERTEXT_WIDTH'd14370606;
publickey_row[1527] = `CIPHERTEXT_WIDTH'd10614891;
publickey_row[1528] = `CIPHERTEXT_WIDTH'd3493727;
publickey_row[1529] = `CIPHERTEXT_WIDTH'd9251468;
publickey_row[1530] = `CIPHERTEXT_WIDTH'd14697209;
publickey_row[1531] = `CIPHERTEXT_WIDTH'd12989616;
publickey_row[1532] = `CIPHERTEXT_WIDTH'd8838881;
publickey_row[1533] = `CIPHERTEXT_WIDTH'd1567072;
publickey_row[1534] = `CIPHERTEXT_WIDTH'd2920908;
publickey_row[1535] = `CIPHERTEXT_WIDTH'd6306933;
publickey_row[1536] = `CIPHERTEXT_WIDTH'd11459002;
publickey_row[1537] = `CIPHERTEXT_WIDTH'd15938927;
publickey_row[1538] = `CIPHERTEXT_WIDTH'd15969139;
publickey_row[1539] = `CIPHERTEXT_WIDTH'd12717796;
publickey_row[1540] = `CIPHERTEXT_WIDTH'd9584073;
publickey_row[1541] = `CIPHERTEXT_WIDTH'd14322869;
publickey_row[1542] = `CIPHERTEXT_WIDTH'd5366833;
publickey_row[1543] = `CIPHERTEXT_WIDTH'd3628330;
publickey_row[1544] = `CIPHERTEXT_WIDTH'd12087565;
publickey_row[1545] = `CIPHERTEXT_WIDTH'd4965187;
publickey_row[1546] = `CIPHERTEXT_WIDTH'd8915878;
publickey_row[1547] = `CIPHERTEXT_WIDTH'd759027;
publickey_row[1548] = `CIPHERTEXT_WIDTH'd2134569;
publickey_row[1549] = `CIPHERTEXT_WIDTH'd2433242;
publickey_row[1550] = `CIPHERTEXT_WIDTH'd16101969;
publickey_row[1551] = `CIPHERTEXT_WIDTH'd5306419;
publickey_row[1552] = `CIPHERTEXT_WIDTH'd8314749;
publickey_row[1553] = `CIPHERTEXT_WIDTH'd2986031;
publickey_row[1554] = `CIPHERTEXT_WIDTH'd5118901;
publickey_row[1555] = `CIPHERTEXT_WIDTH'd14715941;
publickey_row[1556] = `CIPHERTEXT_WIDTH'd9675654;
publickey_row[1557] = `CIPHERTEXT_WIDTH'd15955606;
publickey_row[1558] = `CIPHERTEXT_WIDTH'd4260555;
publickey_row[1559] = `CIPHERTEXT_WIDTH'd6600226;
publickey_row[1560] = `CIPHERTEXT_WIDTH'd14332452;
publickey_row[1561] = `CIPHERTEXT_WIDTH'd4724186;
publickey_row[1562] = `CIPHERTEXT_WIDTH'd14054414;
publickey_row[1563] = `CIPHERTEXT_WIDTH'd5316981;
publickey_row[1564] = `CIPHERTEXT_WIDTH'd9675650;
publickey_row[1565] = `CIPHERTEXT_WIDTH'd8156883;
publickey_row[1566] = `CIPHERTEXT_WIDTH'd8436066;
publickey_row[1567] = `CIPHERTEXT_WIDTH'd2299614;
publickey_row[1568] = `CIPHERTEXT_WIDTH'd2577305;
publickey_row[1569] = `CIPHERTEXT_WIDTH'd16677666;
publickey_row[1570] = `CIPHERTEXT_WIDTH'd15143844;
publickey_row[1571] = `CIPHERTEXT_WIDTH'd5950862;
publickey_row[1572] = `CIPHERTEXT_WIDTH'd7910205;
publickey_row[1573] = `CIPHERTEXT_WIDTH'd945550;
publickey_row[1574] = `CIPHERTEXT_WIDTH'd8659758;
publickey_row[1575] = `CIPHERTEXT_WIDTH'd5236843;
publickey_row[1576] = `CIPHERTEXT_WIDTH'd13784574;
publickey_row[1577] = `CIPHERTEXT_WIDTH'd2575857;
publickey_row[1578] = `CIPHERTEXT_WIDTH'd2117762;
publickey_row[1579] = `CIPHERTEXT_WIDTH'd7398249;
publickey_row[1580] = `CIPHERTEXT_WIDTH'd3780551;
publickey_row[1581] = `CIPHERTEXT_WIDTH'd10458029;
publickey_row[1582] = `CIPHERTEXT_WIDTH'd16402837;
publickey_row[1583] = `CIPHERTEXT_WIDTH'd6616362;
publickey_row[1584] = `CIPHERTEXT_WIDTH'd12053141;
publickey_row[1585] = `CIPHERTEXT_WIDTH'd16219249;
publickey_row[1586] = `CIPHERTEXT_WIDTH'd1399082;
publickey_row[1587] = `CIPHERTEXT_WIDTH'd10599754;
publickey_row[1588] = `CIPHERTEXT_WIDTH'd9207358;
publickey_row[1589] = `CIPHERTEXT_WIDTH'd3762561;
publickey_row[1590] = `CIPHERTEXT_WIDTH'd7610279;
publickey_row[1591] = `CIPHERTEXT_WIDTH'd8155484;
publickey_row[1592] = `CIPHERTEXT_WIDTH'd11675992;
publickey_row[1593] = `CIPHERTEXT_WIDTH'd612512;
publickey_row[1594] = `CIPHERTEXT_WIDTH'd7006755;
publickey_row[1595] = `CIPHERTEXT_WIDTH'd15804566;
publickey_row[1596] = `CIPHERTEXT_WIDTH'd5389904;
publickey_row[1597] = `CIPHERTEXT_WIDTH'd10142299;
publickey_row[1598] = `CIPHERTEXT_WIDTH'd15291721;
publickey_row[1599] = `CIPHERTEXT_WIDTH'd509876;
publickey_row[1600] = `CIPHERTEXT_WIDTH'd10314546;
publickey_row[1601] = `CIPHERTEXT_WIDTH'd13046816;
publickey_row[1602] = `CIPHERTEXT_WIDTH'd15258763;
publickey_row[1603] = `CIPHERTEXT_WIDTH'd14383591;
publickey_row[1604] = `CIPHERTEXT_WIDTH'd16475349;
publickey_row[1605] = `CIPHERTEXT_WIDTH'd11910617;
publickey_row[1606] = `CIPHERTEXT_WIDTH'd8003123;
publickey_row[1607] = `CIPHERTEXT_WIDTH'd14742608;
publickey_row[1608] = `CIPHERTEXT_WIDTH'd4783189;
publickey_row[1609] = `CIPHERTEXT_WIDTH'd7902002;
publickey_row[1610] = `CIPHERTEXT_WIDTH'd3248176;
publickey_row[1611] = `CIPHERTEXT_WIDTH'd8134601;
publickey_row[1612] = `CIPHERTEXT_WIDTH'd845499;
publickey_row[1613] = `CIPHERTEXT_WIDTH'd4867743;
publickey_row[1614] = `CIPHERTEXT_WIDTH'd3703089;
publickey_row[1615] = `CIPHERTEXT_WIDTH'd15437356;
publickey_row[1616] = `CIPHERTEXT_WIDTH'd4936773;
publickey_row[1617] = `CIPHERTEXT_WIDTH'd6734161;
publickey_row[1618] = `CIPHERTEXT_WIDTH'd5175828;
publickey_row[1619] = `CIPHERTEXT_WIDTH'd4327365;
publickey_row[1620] = `CIPHERTEXT_WIDTH'd12828166;
publickey_row[1621] = `CIPHERTEXT_WIDTH'd9614036;
publickey_row[1622] = `CIPHERTEXT_WIDTH'd15089794;
publickey_row[1623] = `CIPHERTEXT_WIDTH'd4295989;
publickey_row[1624] = `CIPHERTEXT_WIDTH'd10711156;
publickey_row[1625] = `CIPHERTEXT_WIDTH'd1046252;
publickey_row[1626] = `CIPHERTEXT_WIDTH'd3149932;
publickey_row[1627] = `CIPHERTEXT_WIDTH'd9738531;
publickey_row[1628] = `CIPHERTEXT_WIDTH'd15104852;
publickey_row[1629] = `CIPHERTEXT_WIDTH'd13897023;
publickey_row[1630] = `CIPHERTEXT_WIDTH'd5163971;
publickey_row[1631] = `CIPHERTEXT_WIDTH'd10647497;
publickey_row[1632] = `CIPHERTEXT_WIDTH'd4930571;
publickey_row[1633] = `CIPHERTEXT_WIDTH'd5093076;
publickey_row[1634] = `CIPHERTEXT_WIDTH'd8237497;
publickey_row[1635] = `CIPHERTEXT_WIDTH'd4837059;
publickey_row[1636] = `CIPHERTEXT_WIDTH'd11722471;
publickey_row[1637] = `CIPHERTEXT_WIDTH'd10836541;
publickey_row[1638] = `CIPHERTEXT_WIDTH'd12084914;
publickey_row[1639] = `CIPHERTEXT_WIDTH'd6670774;
publickey_row[1640] = `CIPHERTEXT_WIDTH'd4151381;
publickey_row[1641] = `CIPHERTEXT_WIDTH'd13549890;
publickey_row[1642] = `CIPHERTEXT_WIDTH'd12719770;
publickey_row[1643] = `CIPHERTEXT_WIDTH'd16357094;
publickey_row[1644] = `CIPHERTEXT_WIDTH'd7814814;
publickey_row[1645] = `CIPHERTEXT_WIDTH'd3667306;
publickey_row[1646] = `CIPHERTEXT_WIDTH'd284332;
publickey_row[1647] = `CIPHERTEXT_WIDTH'd3914720;
publickey_row[1648] = `CIPHERTEXT_WIDTH'd12210385;
publickey_row[1649] = `CIPHERTEXT_WIDTH'd14184284;
publickey_row[1650] = `CIPHERTEXT_WIDTH'd3828168;
publickey_row[1651] = `CIPHERTEXT_WIDTH'd7804221;
publickey_row[1652] = `CIPHERTEXT_WIDTH'd6366040;
publickey_row[1653] = `CIPHERTEXT_WIDTH'd7856735;
publickey_row[1654] = `CIPHERTEXT_WIDTH'd12739530;
publickey_row[1655] = `CIPHERTEXT_WIDTH'd7774134;
publickey_row[1656] = `CIPHERTEXT_WIDTH'd4485613;
publickey_row[1657] = `CIPHERTEXT_WIDTH'd4371191;
publickey_row[1658] = `CIPHERTEXT_WIDTH'd6812689;
publickey_row[1659] = `CIPHERTEXT_WIDTH'd12466371;
publickey_row[1660] = `CIPHERTEXT_WIDTH'd2249828;
publickey_row[1661] = `CIPHERTEXT_WIDTH'd14844870;
publickey_row[1662] = `CIPHERTEXT_WIDTH'd5374584;
publickey_row[1663] = `CIPHERTEXT_WIDTH'd5529359;
publickey_row[1664] = `CIPHERTEXT_WIDTH'd15433273;
publickey_row[1665] = `CIPHERTEXT_WIDTH'd1361806;
publickey_row[1666] = `CIPHERTEXT_WIDTH'd11370001;
publickey_row[1667] = `CIPHERTEXT_WIDTH'd12726994;
publickey_row[1668] = `CIPHERTEXT_WIDTH'd7308420;
publickey_row[1669] = `CIPHERTEXT_WIDTH'd9498106;
publickey_row[1670] = `CIPHERTEXT_WIDTH'd2260172;
publickey_row[1671] = `CIPHERTEXT_WIDTH'd15729047;
publickey_row[1672] = `CIPHERTEXT_WIDTH'd8683997;
publickey_row[1673] = `CIPHERTEXT_WIDTH'd15887361;
publickey_row[1674] = `CIPHERTEXT_WIDTH'd12667794;
publickey_row[1675] = `CIPHERTEXT_WIDTH'd244435;
publickey_row[1676] = `CIPHERTEXT_WIDTH'd14967887;
publickey_row[1677] = `CIPHERTEXT_WIDTH'd4299294;
publickey_row[1678] = `CIPHERTEXT_WIDTH'd6822358;
publickey_row[1679] = `CIPHERTEXT_WIDTH'd2287711;
publickey_row[1680] = `CIPHERTEXT_WIDTH'd15998348;
publickey_row[1681] = `CIPHERTEXT_WIDTH'd5717148;
publickey_row[1682] = `CIPHERTEXT_WIDTH'd15663842;
publickey_row[1683] = `CIPHERTEXT_WIDTH'd2974134;
publickey_row[1684] = `CIPHERTEXT_WIDTH'd5574379;
publickey_row[1685] = `CIPHERTEXT_WIDTH'd4334619;
publickey_row[1686] = `CIPHERTEXT_WIDTH'd13140812;
publickey_row[1687] = `CIPHERTEXT_WIDTH'd8479703;
publickey_row[1688] = `CIPHERTEXT_WIDTH'd11271172;
publickey_row[1689] = `CIPHERTEXT_WIDTH'd15290983;
publickey_row[1690] = `CIPHERTEXT_WIDTH'd1305759;
publickey_row[1691] = `CIPHERTEXT_WIDTH'd13701625;
publickey_row[1692] = `CIPHERTEXT_WIDTH'd14274269;
publickey_row[1693] = `CIPHERTEXT_WIDTH'd6661629;
publickey_row[1694] = `CIPHERTEXT_WIDTH'd8542544;
publickey_row[1695] = `CIPHERTEXT_WIDTH'd15471564;
publickey_row[1696] = `CIPHERTEXT_WIDTH'd11643863;
publickey_row[1697] = `CIPHERTEXT_WIDTH'd8444283;
publickey_row[1698] = `CIPHERTEXT_WIDTH'd2180914;
publickey_row[1699] = `CIPHERTEXT_WIDTH'd9631593;
publickey_row[1700] = `CIPHERTEXT_WIDTH'd9693412;
publickey_row[1701] = `CIPHERTEXT_WIDTH'd4913701;
publickey_row[1702] = `CIPHERTEXT_WIDTH'd12880978;
publickey_row[1703] = `CIPHERTEXT_WIDTH'd14888923;
publickey_row[1704] = `CIPHERTEXT_WIDTH'd8301348;
publickey_row[1705] = `CIPHERTEXT_WIDTH'd13418293;
publickey_row[1706] = `CIPHERTEXT_WIDTH'd5869934;
publickey_row[1707] = `CIPHERTEXT_WIDTH'd12257776;
publickey_row[1708] = `CIPHERTEXT_WIDTH'd13761273;
publickey_row[1709] = `CIPHERTEXT_WIDTH'd5773742;
publickey_row[1710] = `CIPHERTEXT_WIDTH'd14284263;
publickey_row[1711] = `CIPHERTEXT_WIDTH'd14632099;
publickey_row[1712] = `CIPHERTEXT_WIDTH'd5008389;
publickey_row[1713] = `CIPHERTEXT_WIDTH'd1575479;
publickey_row[1714] = `CIPHERTEXT_WIDTH'd8425394;
publickey_row[1715] = `CIPHERTEXT_WIDTH'd7807855;
publickey_row[1716] = `CIPHERTEXT_WIDTH'd10916233;
publickey_row[1717] = `CIPHERTEXT_WIDTH'd12775755;
publickey_row[1718] = `CIPHERTEXT_WIDTH'd16542474;
publickey_row[1719] = `CIPHERTEXT_WIDTH'd6779875;
publickey_row[1720] = `CIPHERTEXT_WIDTH'd16290959;
publickey_row[1721] = `CIPHERTEXT_WIDTH'd16722605;
publickey_row[1722] = `CIPHERTEXT_WIDTH'd11745459;
publickey_row[1723] = `CIPHERTEXT_WIDTH'd11350808;
publickey_row[1724] = `CIPHERTEXT_WIDTH'd158732;
publickey_row[1725] = `CIPHERTEXT_WIDTH'd5522075;
publickey_row[1726] = `CIPHERTEXT_WIDTH'd4891201;
publickey_row[1727] = `CIPHERTEXT_WIDTH'd10900772;
publickey_row[1728] = `CIPHERTEXT_WIDTH'd2680330;
publickey_row[1729] = `CIPHERTEXT_WIDTH'd7206193;
publickey_row[1730] = `CIPHERTEXT_WIDTH'd15659914;
publickey_row[1731] = `CIPHERTEXT_WIDTH'd2875614;
publickey_row[1732] = `CIPHERTEXT_WIDTH'd13546980;
publickey_row[1733] = `CIPHERTEXT_WIDTH'd2974732;
publickey_row[1734] = `CIPHERTEXT_WIDTH'd1582435;
publickey_row[1735] = `CIPHERTEXT_WIDTH'd16289363;
publickey_row[1736] = `CIPHERTEXT_WIDTH'd9155741;
publickey_row[1737] = `CIPHERTEXT_WIDTH'd9734084;
publickey_row[1738] = `CIPHERTEXT_WIDTH'd6552390;
publickey_row[1739] = `CIPHERTEXT_WIDTH'd7665480;
publickey_row[1740] = `CIPHERTEXT_WIDTH'd1564433;
publickey_row[1741] = `CIPHERTEXT_WIDTH'd6466971;
publickey_row[1742] = `CIPHERTEXT_WIDTH'd12855230;
publickey_row[1743] = `CIPHERTEXT_WIDTH'd14136634;
publickey_row[1744] = `CIPHERTEXT_WIDTH'd12063251;
publickey_row[1745] = `CIPHERTEXT_WIDTH'd9322549;
publickey_row[1746] = `CIPHERTEXT_WIDTH'd5514083;
publickey_row[1747] = `CIPHERTEXT_WIDTH'd13323338;
publickey_row[1748] = `CIPHERTEXT_WIDTH'd2905902;
publickey_row[1749] = `CIPHERTEXT_WIDTH'd6971800;
publickey_row[1750] = `CIPHERTEXT_WIDTH'd5500325;
publickey_row[1751] = `CIPHERTEXT_WIDTH'd1804103;
publickey_row[1752] = `CIPHERTEXT_WIDTH'd2028603;
publickey_row[1753] = `CIPHERTEXT_WIDTH'd9934175;
publickey_row[1754] = `CIPHERTEXT_WIDTH'd6395941;
publickey_row[1755] = `CIPHERTEXT_WIDTH'd13045594;
publickey_row[1756] = `CIPHERTEXT_WIDTH'd5507242;
publickey_row[1757] = `CIPHERTEXT_WIDTH'd2357792;
publickey_row[1758] = `CIPHERTEXT_WIDTH'd14761477;
publickey_row[1759] = `CIPHERTEXT_WIDTH'd9323467;
publickey_row[1760] = `CIPHERTEXT_WIDTH'd858965;
publickey_row[1761] = `CIPHERTEXT_WIDTH'd7356477;
publickey_row[1762] = `CIPHERTEXT_WIDTH'd14028938;
publickey_row[1763] = `CIPHERTEXT_WIDTH'd8725112;
publickey_row[1764] = `CIPHERTEXT_WIDTH'd14112192;
publickey_row[1765] = `CIPHERTEXT_WIDTH'd4759116;
publickey_row[1766] = `CIPHERTEXT_WIDTH'd10562941;
publickey_row[1767] = `CIPHERTEXT_WIDTH'd9402381;
publickey_row[1768] = `CIPHERTEXT_WIDTH'd1109328;
publickey_row[1769] = `CIPHERTEXT_WIDTH'd7952783;
publickey_row[1770] = `CIPHERTEXT_WIDTH'd1987673;
publickey_row[1771] = `CIPHERTEXT_WIDTH'd6215640;
publickey_row[1772] = `CIPHERTEXT_WIDTH'd15332430;
publickey_row[1773] = `CIPHERTEXT_WIDTH'd12148586;
publickey_row[1774] = `CIPHERTEXT_WIDTH'd8618655;
publickey_row[1775] = `CIPHERTEXT_WIDTH'd7540392;
publickey_row[1776] = `CIPHERTEXT_WIDTH'd13072315;
publickey_row[1777] = `CIPHERTEXT_WIDTH'd13110044;
publickey_row[1778] = `CIPHERTEXT_WIDTH'd14125567;
publickey_row[1779] = `CIPHERTEXT_WIDTH'd8362306;
publickey_row[1780] = `CIPHERTEXT_WIDTH'd10268540;
publickey_row[1781] = `CIPHERTEXT_WIDTH'd973922;
publickey_row[1782] = `CIPHERTEXT_WIDTH'd7809937;
publickey_row[1783] = `CIPHERTEXT_WIDTH'd10199032;
publickey_row[1784] = `CIPHERTEXT_WIDTH'd8564653;
publickey_row[1785] = `CIPHERTEXT_WIDTH'd4495821;
publickey_row[1786] = `CIPHERTEXT_WIDTH'd4661668;
publickey_row[1787] = `CIPHERTEXT_WIDTH'd11581870;
publickey_row[1788] = `CIPHERTEXT_WIDTH'd2633309;
publickey_row[1789] = `CIPHERTEXT_WIDTH'd4706862;
publickey_row[1790] = `CIPHERTEXT_WIDTH'd11910366;
publickey_row[1791] = `CIPHERTEXT_WIDTH'd8985979;
publickey_row[1792] = `CIPHERTEXT_WIDTH'd6195224;
publickey_row[1793] = `CIPHERTEXT_WIDTH'd2888608;
publickey_row[1794] = `CIPHERTEXT_WIDTH'd6929444;
publickey_row[1795] = `CIPHERTEXT_WIDTH'd3324596;
publickey_row[1796] = `CIPHERTEXT_WIDTH'd6533180;
publickey_row[1797] = `CIPHERTEXT_WIDTH'd12344974;
publickey_row[1798] = `CIPHERTEXT_WIDTH'd2700443;
publickey_row[1799] = `CIPHERTEXT_WIDTH'd11862733;
publickey_row[1800] = `CIPHERTEXT_WIDTH'd13551769;
publickey_row[1801] = `CIPHERTEXT_WIDTH'd12856810;
publickey_row[1802] = `CIPHERTEXT_WIDTH'd3665952;
publickey_row[1803] = `CIPHERTEXT_WIDTH'd4887133;
publickey_row[1804] = `CIPHERTEXT_WIDTH'd4607618;
publickey_row[1805] = `CIPHERTEXT_WIDTH'd15147691;
publickey_row[1806] = `CIPHERTEXT_WIDTH'd3126521;
publickey_row[1807] = `CIPHERTEXT_WIDTH'd10569500;
publickey_row[1808] = `CIPHERTEXT_WIDTH'd632842;
publickey_row[1809] = `CIPHERTEXT_WIDTH'd3539842;
publickey_row[1810] = `CIPHERTEXT_WIDTH'd13468313;
publickey_row[1811] = `CIPHERTEXT_WIDTH'd15341379;
publickey_row[1812] = `CIPHERTEXT_WIDTH'd6568976;
publickey_row[1813] = `CIPHERTEXT_WIDTH'd3942788;
publickey_row[1814] = `CIPHERTEXT_WIDTH'd14462304;
publickey_row[1815] = `CIPHERTEXT_WIDTH'd1628205;
publickey_row[1816] = `CIPHERTEXT_WIDTH'd6267558;
publickey_row[1817] = `CIPHERTEXT_WIDTH'd10887295;
publickey_row[1818] = `CIPHERTEXT_WIDTH'd14676162;
publickey_row[1819] = `CIPHERTEXT_WIDTH'd2222093;
publickey_row[1820] = `CIPHERTEXT_WIDTH'd12748329;
publickey_row[1821] = `CIPHERTEXT_WIDTH'd1321065;
publickey_row[1822] = `CIPHERTEXT_WIDTH'd3912072;
publickey_row[1823] = `CIPHERTEXT_WIDTH'd9263274;
publickey_row[1824] = `CIPHERTEXT_WIDTH'd12075058;
publickey_row[1825] = `CIPHERTEXT_WIDTH'd10974709;
publickey_row[1826] = `CIPHERTEXT_WIDTH'd9496843;
publickey_row[1827] = `CIPHERTEXT_WIDTH'd7859566;
publickey_row[1828] = `CIPHERTEXT_WIDTH'd8693097;
publickey_row[1829] = `CIPHERTEXT_WIDTH'd3519897;
publickey_row[1830] = `CIPHERTEXT_WIDTH'd14512064;
publickey_row[1831] = `CIPHERTEXT_WIDTH'd16191947;
publickey_row[1832] = `CIPHERTEXT_WIDTH'd1695851;
publickey_row[1833] = `CIPHERTEXT_WIDTH'd3233092;
publickey_row[1834] = `CIPHERTEXT_WIDTH'd1570307;
publickey_row[1835] = `CIPHERTEXT_WIDTH'd12073701;
publickey_row[1836] = `CIPHERTEXT_WIDTH'd5429874;
publickey_row[1837] = `CIPHERTEXT_WIDTH'd311753;
publickey_row[1838] = `CIPHERTEXT_WIDTH'd12055720;
publickey_row[1839] = `CIPHERTEXT_WIDTH'd12437439;
publickey_row[1840] = `CIPHERTEXT_WIDTH'd2808672;
publickey_row[1841] = `CIPHERTEXT_WIDTH'd6439803;
publickey_row[1842] = `CIPHERTEXT_WIDTH'd15983986;
publickey_row[1843] = `CIPHERTEXT_WIDTH'd2847381;
publickey_row[1844] = `CIPHERTEXT_WIDTH'd9381697;
publickey_row[1845] = `CIPHERTEXT_WIDTH'd11968172;
publickey_row[1846] = `CIPHERTEXT_WIDTH'd16181977;
publickey_row[1847] = `CIPHERTEXT_WIDTH'd8948253;
publickey_row[1848] = `CIPHERTEXT_WIDTH'd15446586;
publickey_row[1849] = `CIPHERTEXT_WIDTH'd5074562;
publickey_row[1850] = `CIPHERTEXT_WIDTH'd1304363;
publickey_row[1851] = `CIPHERTEXT_WIDTH'd14751308;
publickey_row[1852] = `CIPHERTEXT_WIDTH'd15964611;
publickey_row[1853] = `CIPHERTEXT_WIDTH'd12375585;
publickey_row[1854] = `CIPHERTEXT_WIDTH'd10708275;
publickey_row[1855] = `CIPHERTEXT_WIDTH'd3447692;
publickey_row[1856] = `CIPHERTEXT_WIDTH'd9339147;
publickey_row[1857] = `CIPHERTEXT_WIDTH'd3474867;
publickey_row[1858] = `CIPHERTEXT_WIDTH'd3601629;
publickey_row[1859] = `CIPHERTEXT_WIDTH'd4355453;
publickey_row[1860] = `CIPHERTEXT_WIDTH'd13447058;
publickey_row[1861] = `CIPHERTEXT_WIDTH'd15774664;
publickey_row[1862] = `CIPHERTEXT_WIDTH'd6877265;
publickey_row[1863] = `CIPHERTEXT_WIDTH'd7510546;
publickey_row[1864] = `CIPHERTEXT_WIDTH'd10854773;
publickey_row[1865] = `CIPHERTEXT_WIDTH'd14235787;
publickey_row[1866] = `CIPHERTEXT_WIDTH'd7554646;
publickey_row[1867] = `CIPHERTEXT_WIDTH'd13327660;
publickey_row[1868] = `CIPHERTEXT_WIDTH'd13689138;
publickey_row[1869] = `CIPHERTEXT_WIDTH'd14506554;
publickey_row[1870] = `CIPHERTEXT_WIDTH'd344899;
publickey_row[1871] = `CIPHERTEXT_WIDTH'd5719583;
publickey_row[1872] = `CIPHERTEXT_WIDTH'd1272825;
publickey_row[1873] = `CIPHERTEXT_WIDTH'd11852713;
publickey_row[1874] = `CIPHERTEXT_WIDTH'd758793;
publickey_row[1875] = `CIPHERTEXT_WIDTH'd9376385;
publickey_row[1876] = `CIPHERTEXT_WIDTH'd8176268;
publickey_row[1877] = `CIPHERTEXT_WIDTH'd10623835;
publickey_row[1878] = `CIPHERTEXT_WIDTH'd8218194;
publickey_row[1879] = `CIPHERTEXT_WIDTH'd11966204;
publickey_row[1880] = `CIPHERTEXT_WIDTH'd8426163;
publickey_row[1881] = `CIPHERTEXT_WIDTH'd7310930;
publickey_row[1882] = `CIPHERTEXT_WIDTH'd3469316;
publickey_row[1883] = `CIPHERTEXT_WIDTH'd313998;
publickey_row[1884] = `CIPHERTEXT_WIDTH'd5207567;
publickey_row[1885] = `CIPHERTEXT_WIDTH'd2076398;
publickey_row[1886] = `CIPHERTEXT_WIDTH'd11945763;
publickey_row[1887] = `CIPHERTEXT_WIDTH'd12355957;
publickey_row[1888] = `CIPHERTEXT_WIDTH'd11131683;
publickey_row[1889] = `CIPHERTEXT_WIDTH'd8234898;
publickey_row[1890] = `CIPHERTEXT_WIDTH'd13818856;
publickey_row[1891] = `CIPHERTEXT_WIDTH'd1231155;
publickey_row[1892] = `CIPHERTEXT_WIDTH'd6273303;
publickey_row[1893] = `CIPHERTEXT_WIDTH'd16769458;
publickey_row[1894] = `CIPHERTEXT_WIDTH'd798779;
publickey_row[1895] = `CIPHERTEXT_WIDTH'd14742223;
publickey_row[1896] = `CIPHERTEXT_WIDTH'd16315110;
publickey_row[1897] = `CIPHERTEXT_WIDTH'd2167783;
publickey_row[1898] = `CIPHERTEXT_WIDTH'd7102901;
publickey_row[1899] = `CIPHERTEXT_WIDTH'd11878841;
publickey_row[1900] = `CIPHERTEXT_WIDTH'd10283012;
publickey_row[1901] = `CIPHERTEXT_WIDTH'd10624609;
publickey_row[1902] = `CIPHERTEXT_WIDTH'd13165656;
publickey_row[1903] = `CIPHERTEXT_WIDTH'd16507595;
publickey_row[1904] = `CIPHERTEXT_WIDTH'd15777198;
publickey_row[1905] = `CIPHERTEXT_WIDTH'd15881358;
publickey_row[1906] = `CIPHERTEXT_WIDTH'd9399046;
publickey_row[1907] = `CIPHERTEXT_WIDTH'd12011940;
publickey_row[1908] = `CIPHERTEXT_WIDTH'd13241141;
publickey_row[1909] = `CIPHERTEXT_WIDTH'd8004562;
publickey_row[1910] = `CIPHERTEXT_WIDTH'd16717516;
publickey_row[1911] = `CIPHERTEXT_WIDTH'd12823941;
publickey_row[1912] = `CIPHERTEXT_WIDTH'd4711942;
publickey_row[1913] = `CIPHERTEXT_WIDTH'd9067364;
publickey_row[1914] = `CIPHERTEXT_WIDTH'd11197599;
publickey_row[1915] = `CIPHERTEXT_WIDTH'd7509891;
publickey_row[1916] = `CIPHERTEXT_WIDTH'd15127635;
publickey_row[1917] = `CIPHERTEXT_WIDTH'd14373282;
publickey_row[1918] = `CIPHERTEXT_WIDTH'd8933307;
publickey_row[1919] = `CIPHERTEXT_WIDTH'd5323359;
publickey_row[1920] = `CIPHERTEXT_WIDTH'd13043164;
publickey_row[1921] = `CIPHERTEXT_WIDTH'd9551435;
publickey_row[1922] = `CIPHERTEXT_WIDTH'd6394494;
publickey_row[1923] = `CIPHERTEXT_WIDTH'd15141845;
publickey_row[1924] = `CIPHERTEXT_WIDTH'd173633;
publickey_row[1925] = `CIPHERTEXT_WIDTH'd12662654;
publickey_row[1926] = `CIPHERTEXT_WIDTH'd14376281;
publickey_row[1927] = `CIPHERTEXT_WIDTH'd2254940;
publickey_row[1928] = `CIPHERTEXT_WIDTH'd2009592;
publickey_row[1929] = `CIPHERTEXT_WIDTH'd12593908;
publickey_row[1930] = `CIPHERTEXT_WIDTH'd1768107;
publickey_row[1931] = `CIPHERTEXT_WIDTH'd7568063;
publickey_row[1932] = `CIPHERTEXT_WIDTH'd11936452;
publickey_row[1933] = `CIPHERTEXT_WIDTH'd10905349;
publickey_row[1934] = `CIPHERTEXT_WIDTH'd13517104;
publickey_row[1935] = `CIPHERTEXT_WIDTH'd948922;
publickey_row[1936] = `CIPHERTEXT_WIDTH'd794864;
publickey_row[1937] = `CIPHERTEXT_WIDTH'd160131;
publickey_row[1938] = `CIPHERTEXT_WIDTH'd4560735;
publickey_row[1939] = `CIPHERTEXT_WIDTH'd1673228;
publickey_row[1940] = `CIPHERTEXT_WIDTH'd7001501;
publickey_row[1941] = `CIPHERTEXT_WIDTH'd3496702;
publickey_row[1942] = `CIPHERTEXT_WIDTH'd4285683;
publickey_row[1943] = `CIPHERTEXT_WIDTH'd563333;
publickey_row[1944] = `CIPHERTEXT_WIDTH'd10966394;
publickey_row[1945] = `CIPHERTEXT_WIDTH'd16366651;
publickey_row[1946] = `CIPHERTEXT_WIDTH'd533638;
publickey_row[1947] = `CIPHERTEXT_WIDTH'd2143402;
publickey_row[1948] = `CIPHERTEXT_WIDTH'd10770434;
publickey_row[1949] = `CIPHERTEXT_WIDTH'd12767296;
publickey_row[1950] = `CIPHERTEXT_WIDTH'd10771265;
publickey_row[1951] = `CIPHERTEXT_WIDTH'd14233564;
publickey_row[1952] = `CIPHERTEXT_WIDTH'd11360186;
publickey_row[1953] = `CIPHERTEXT_WIDTH'd5973164;
publickey_row[1954] = `CIPHERTEXT_WIDTH'd6979749;
publickey_row[1955] = `CIPHERTEXT_WIDTH'd1881130;
publickey_row[1956] = `CIPHERTEXT_WIDTH'd10334923;
publickey_row[1957] = `CIPHERTEXT_WIDTH'd7744809;
publickey_row[1958] = `CIPHERTEXT_WIDTH'd680315;
publickey_row[1959] = `CIPHERTEXT_WIDTH'd12964780;
publickey_row[1960] = `CIPHERTEXT_WIDTH'd9570480;
publickey_row[1961] = `CIPHERTEXT_WIDTH'd15419914;
publickey_row[1962] = `CIPHERTEXT_WIDTH'd3459339;
publickey_row[1963] = `CIPHERTEXT_WIDTH'd8028590;
publickey_row[1964] = `CIPHERTEXT_WIDTH'd4050903;
publickey_row[1965] = `CIPHERTEXT_WIDTH'd15058069;
publickey_row[1966] = `CIPHERTEXT_WIDTH'd1490641;
publickey_row[1967] = `CIPHERTEXT_WIDTH'd5425825;
publickey_row[1968] = `CIPHERTEXT_WIDTH'd12465754;
publickey_row[1969] = `CIPHERTEXT_WIDTH'd2215942;
publickey_row[1970] = `CIPHERTEXT_WIDTH'd7953107;
publickey_row[1971] = `CIPHERTEXT_WIDTH'd2649305;
publickey_row[1972] = `CIPHERTEXT_WIDTH'd12219061;
publickey_row[1973] = `CIPHERTEXT_WIDTH'd15247206;
publickey_row[1974] = `CIPHERTEXT_WIDTH'd13517978;
publickey_row[1975] = `CIPHERTEXT_WIDTH'd10033135;
publickey_row[1976] = `CIPHERTEXT_WIDTH'd1356883;
publickey_row[1977] = `CIPHERTEXT_WIDTH'd13334495;
publickey_row[1978] = `CIPHERTEXT_WIDTH'd13071694;
publickey_row[1979] = `CIPHERTEXT_WIDTH'd12163158;
publickey_row[1980] = `CIPHERTEXT_WIDTH'd15965064;
publickey_row[1981] = `CIPHERTEXT_WIDTH'd6892900;
publickey_row[1982] = `CIPHERTEXT_WIDTH'd5460286;
publickey_row[1983] = `CIPHERTEXT_WIDTH'd244826;
publickey_row[1984] = `CIPHERTEXT_WIDTH'd15996325;
publickey_row[1985] = `CIPHERTEXT_WIDTH'd12273083;
publickey_row[1986] = `CIPHERTEXT_WIDTH'd2276601;
publickey_row[1987] = `CIPHERTEXT_WIDTH'd273011;
publickey_row[1988] = `CIPHERTEXT_WIDTH'd3683288;
publickey_row[1989] = `CIPHERTEXT_WIDTH'd3124026;
publickey_row[1990] = `CIPHERTEXT_WIDTH'd11258733;
publickey_row[1991] = `CIPHERTEXT_WIDTH'd9322656;
publickey_row[1992] = `CIPHERTEXT_WIDTH'd2917605;
publickey_row[1993] = `CIPHERTEXT_WIDTH'd9056899;
publickey_row[1994] = `CIPHERTEXT_WIDTH'd5252203;
publickey_row[1995] = `CIPHERTEXT_WIDTH'd10282608;
publickey_row[1996] = `CIPHERTEXT_WIDTH'd8217695;
publickey_row[1997] = `CIPHERTEXT_WIDTH'd9451589;
publickey_row[1998] = `CIPHERTEXT_WIDTH'd7774631;
publickey_row[1999] = `CIPHERTEXT_WIDTH'd14210054;
publickey_row[2000] = `CIPHERTEXT_WIDTH'd10100810;
publickey_row[2001] = `CIPHERTEXT_WIDTH'd8683327;
publickey_row[2002] = `CIPHERTEXT_WIDTH'd5083063;
publickey_row[2003] = `CIPHERTEXT_WIDTH'd14089656;
publickey_row[2004] = `CIPHERTEXT_WIDTH'd13958259;
publickey_row[2005] = `CIPHERTEXT_WIDTH'd11957235;
publickey_row[2006] = `CIPHERTEXT_WIDTH'd13667491;
publickey_row[2007] = `CIPHERTEXT_WIDTH'd2614369;
publickey_row[2008] = `CIPHERTEXT_WIDTH'd7045794;
publickey_row[2009] = `CIPHERTEXT_WIDTH'd5209471;
publickey_row[2010] = `CIPHERTEXT_WIDTH'd7365591;
publickey_row[2011] = `CIPHERTEXT_WIDTH'd7621839;
publickey_row[2012] = `CIPHERTEXT_WIDTH'd5738107;
publickey_row[2013] = `CIPHERTEXT_WIDTH'd15527995;
publickey_row[2014] = `CIPHERTEXT_WIDTH'd10523688;
publickey_row[2015] = `CIPHERTEXT_WIDTH'd16169644;
publickey_row[2016] = `CIPHERTEXT_WIDTH'd2136372;
publickey_row[2017] = `CIPHERTEXT_WIDTH'd4095000;
publickey_row[2018] = `CIPHERTEXT_WIDTH'd8236730;
publickey_row[2019] = `CIPHERTEXT_WIDTH'd13122016;
publickey_row[2020] = `CIPHERTEXT_WIDTH'd12278375;
publickey_row[2021] = `CIPHERTEXT_WIDTH'd5411360;
publickey_row[2022] = `CIPHERTEXT_WIDTH'd4415864;
publickey_row[2023] = `CIPHERTEXT_WIDTH'd16308147;
publickey_row[2024] = `CIPHERTEXT_WIDTH'd12250524;
publickey_row[2025] = `CIPHERTEXT_WIDTH'd5775635;
publickey_row[2026] = `CIPHERTEXT_WIDTH'd16003018;
publickey_row[2027] = `CIPHERTEXT_WIDTH'd15857030;
publickey_row[2028] = `CIPHERTEXT_WIDTH'd2733084;
publickey_row[2029] = `CIPHERTEXT_WIDTH'd10161506;
publickey_row[2030] = `CIPHERTEXT_WIDTH'd10747249;
publickey_row[2031] = `CIPHERTEXT_WIDTH'd7077368;
publickey_row[2032] = `CIPHERTEXT_WIDTH'd12125908;
publickey_row[2033] = `CIPHERTEXT_WIDTH'd8522579;
publickey_row[2034] = `CIPHERTEXT_WIDTH'd5734215;
publickey_row[2035] = `CIPHERTEXT_WIDTH'd3720295;
publickey_row[2036] = `CIPHERTEXT_WIDTH'd11527167;
publickey_row[2037] = `CIPHERTEXT_WIDTH'd16014488;
publickey_row[2038] = `CIPHERTEXT_WIDTH'd5249427;
publickey_row[2039] = `CIPHERTEXT_WIDTH'd7091335;
publickey_row[2040] = `CIPHERTEXT_WIDTH'd15467785;
publickey_row[2041] = `CIPHERTEXT_WIDTH'd8459730;
publickey_row[2042] = `CIPHERTEXT_WIDTH'd5155367;
publickey_row[2043] = `CIPHERTEXT_WIDTH'd2914289;
publickey_row[2044] = `CIPHERTEXT_WIDTH'd11735432;
publickey_row[2045] = `CIPHERTEXT_WIDTH'd2935388;
publickey_row[2046] = `CIPHERTEXT_WIDTH'd1878402;
publickey_row[2047] = `CIPHERTEXT_WIDTH'd7240897;
publickey_row[2048] = `CIPHERTEXT_WIDTH'd12616432;
publickey_row[2049] = `CIPHERTEXT_WIDTH'd8999510;
publickey_row[2050] = `CIPHERTEXT_WIDTH'd12702354;
publickey_row[2051] = `CIPHERTEXT_WIDTH'd8290019;
publickey_row[2052] = `CIPHERTEXT_WIDTH'd8958315;
publickey_row[2053] = `CIPHERTEXT_WIDTH'd14667234;
publickey_row[2054] = `CIPHERTEXT_WIDTH'd11335111;
publickey_row[2055] = `CIPHERTEXT_WIDTH'd15994266;
publickey_row[2056] = `CIPHERTEXT_WIDTH'd7151;
publickey_row[2057] = `CIPHERTEXT_WIDTH'd589610;
publickey_row[2058] = `CIPHERTEXT_WIDTH'd9730264;
publickey_row[2059] = `CIPHERTEXT_WIDTH'd10314669;
publickey_row[2060] = `CIPHERTEXT_WIDTH'd3692957;
publickey_row[2061] = `CIPHERTEXT_WIDTH'd7767502;
publickey_row[2062] = `CIPHERTEXT_WIDTH'd11314423;
publickey_row[2063] = `CIPHERTEXT_WIDTH'd1620594;
publickey_row[2064] = `CIPHERTEXT_WIDTH'd15359853;
publickey_row[2065] = `CIPHERTEXT_WIDTH'd3032710;
publickey_row[2066] = `CIPHERTEXT_WIDTH'd1472427;
publickey_row[2067] = `CIPHERTEXT_WIDTH'd11813587;
publickey_row[2068] = `CIPHERTEXT_WIDTH'd7033114;
publickey_row[2069] = `CIPHERTEXT_WIDTH'd15190859;
publickey_row[2070] = `CIPHERTEXT_WIDTH'd8887304;
publickey_row[2071] = `CIPHERTEXT_WIDTH'd12496961;
publickey_row[2072] = `CIPHERTEXT_WIDTH'd10560635;
publickey_row[2073] = `CIPHERTEXT_WIDTH'd6350890;
publickey_row[2074] = `CIPHERTEXT_WIDTH'd16719049;
publickey_row[2075] = `CIPHERTEXT_WIDTH'd10851476;
publickey_row[2076] = `CIPHERTEXT_WIDTH'd15264588;
publickey_row[2077] = `CIPHERTEXT_WIDTH'd6054564;
publickey_row[2078] = `CIPHERTEXT_WIDTH'd8776132;
publickey_row[2079] = `CIPHERTEXT_WIDTH'd1066655;
publickey_row[2080] = `CIPHERTEXT_WIDTH'd13063996;
publickey_row[2081] = `CIPHERTEXT_WIDTH'd306562;
publickey_row[2082] = `CIPHERTEXT_WIDTH'd14876970;
publickey_row[2083] = `CIPHERTEXT_WIDTH'd14188746;
publickey_row[2084] = `CIPHERTEXT_WIDTH'd8615817;
publickey_row[2085] = `CIPHERTEXT_WIDTH'd12438807;
publickey_row[2086] = `CIPHERTEXT_WIDTH'd8443587;
publickey_row[2087] = `CIPHERTEXT_WIDTH'd9714243;
publickey_row[2088] = `CIPHERTEXT_WIDTH'd14015103;
publickey_row[2089] = `CIPHERTEXT_WIDTH'd10466090;
publickey_row[2090] = `CIPHERTEXT_WIDTH'd12024431;
publickey_row[2091] = `CIPHERTEXT_WIDTH'd13042666;
publickey_row[2092] = `CIPHERTEXT_WIDTH'd16247163;
publickey_row[2093] = `CIPHERTEXT_WIDTH'd12600639;
publickey_row[2094] = `CIPHERTEXT_WIDTH'd11853053;
publickey_row[2095] = `CIPHERTEXT_WIDTH'd3337487;
publickey_row[2096] = `CIPHERTEXT_WIDTH'd11004966;
publickey_row[2097] = `CIPHERTEXT_WIDTH'd944201;
publickey_row[2098] = `CIPHERTEXT_WIDTH'd5163542;
publickey_row[2099] = `CIPHERTEXT_WIDTH'd4761469;
publickey_row[2100] = `CIPHERTEXT_WIDTH'd11246777;
publickey_row[2101] = `CIPHERTEXT_WIDTH'd14464162;
publickey_row[2102] = `CIPHERTEXT_WIDTH'd4416222;
publickey_row[2103] = `CIPHERTEXT_WIDTH'd10696380;
publickey_row[2104] = `CIPHERTEXT_WIDTH'd10301180;
publickey_row[2105] = `CIPHERTEXT_WIDTH'd2534191;
publickey_row[2106] = `CIPHERTEXT_WIDTH'd14454704;
publickey_row[2107] = `CIPHERTEXT_WIDTH'd15475653;
publickey_row[2108] = `CIPHERTEXT_WIDTH'd8292014;
publickey_row[2109] = `CIPHERTEXT_WIDTH'd2103166;
publickey_row[2110] = `CIPHERTEXT_WIDTH'd15690991;
publickey_row[2111] = `CIPHERTEXT_WIDTH'd2124566;
publickey_row[2112] = `CIPHERTEXT_WIDTH'd3130437;
publickey_row[2113] = `CIPHERTEXT_WIDTH'd14068734;
publickey_row[2114] = `CIPHERTEXT_WIDTH'd9242399;
publickey_row[2115] = `CIPHERTEXT_WIDTH'd14792110;
publickey_row[2116] = `CIPHERTEXT_WIDTH'd3714020;
publickey_row[2117] = `CIPHERTEXT_WIDTH'd1182739;
publickey_row[2118] = `CIPHERTEXT_WIDTH'd12097281;
publickey_row[2119] = `CIPHERTEXT_WIDTH'd9411381;
publickey_row[2120] = `CIPHERTEXT_WIDTH'd9812960;
publickey_row[2121] = `CIPHERTEXT_WIDTH'd8375635;
publickey_row[2122] = `CIPHERTEXT_WIDTH'd877690;
publickey_row[2123] = `CIPHERTEXT_WIDTH'd8144960;
publickey_row[2124] = `CIPHERTEXT_WIDTH'd5572170;
publickey_row[2125] = `CIPHERTEXT_WIDTH'd8210894;
publickey_row[2126] = `CIPHERTEXT_WIDTH'd6670991;
publickey_row[2127] = `CIPHERTEXT_WIDTH'd46284;
publickey_row[2128] = `CIPHERTEXT_WIDTH'd2614681;
publickey_row[2129] = `CIPHERTEXT_WIDTH'd4026648;
publickey_row[2130] = `CIPHERTEXT_WIDTH'd3602479;
publickey_row[2131] = `CIPHERTEXT_WIDTH'd16142722;
publickey_row[2132] = `CIPHERTEXT_WIDTH'd2847089;
publickey_row[2133] = `CIPHERTEXT_WIDTH'd13800858;
publickey_row[2134] = `CIPHERTEXT_WIDTH'd6657455;
publickey_row[2135] = `CIPHERTEXT_WIDTH'd5615530;
publickey_row[2136] = `CIPHERTEXT_WIDTH'd16035906;
publickey_row[2137] = `CIPHERTEXT_WIDTH'd9119934;
publickey_row[2138] = `CIPHERTEXT_WIDTH'd152859;
publickey_row[2139] = `CIPHERTEXT_WIDTH'd1371282;
publickey_row[2140] = `CIPHERTEXT_WIDTH'd7918821;
publickey_row[2141] = `CIPHERTEXT_WIDTH'd8441930;
publickey_row[2142] = `CIPHERTEXT_WIDTH'd10168998;
publickey_row[2143] = `CIPHERTEXT_WIDTH'd10047465;
publickey_row[2144] = `CIPHERTEXT_WIDTH'd1767100;
publickey_row[2145] = `CIPHERTEXT_WIDTH'd12585545;
publickey_row[2146] = `CIPHERTEXT_WIDTH'd16135636;
publickey_row[2147] = `CIPHERTEXT_WIDTH'd7911838;
publickey_row[2148] = `CIPHERTEXT_WIDTH'd15584299;
publickey_row[2149] = `CIPHERTEXT_WIDTH'd2231317;
publickey_row[2150] = `CIPHERTEXT_WIDTH'd8798799;
publickey_row[2151] = `CIPHERTEXT_WIDTH'd6720404;
publickey_row[2152] = `CIPHERTEXT_WIDTH'd10872142;
publickey_row[2153] = `CIPHERTEXT_WIDTH'd4169323;
publickey_row[2154] = `CIPHERTEXT_WIDTH'd8252980;
publickey_row[2155] = `CIPHERTEXT_WIDTH'd3059133;
publickey_row[2156] = `CIPHERTEXT_WIDTH'd10666849;
publickey_row[2157] = `CIPHERTEXT_WIDTH'd5835831;
publickey_row[2158] = `CIPHERTEXT_WIDTH'd13575720;
publickey_row[2159] = `CIPHERTEXT_WIDTH'd5443121;
publickey_row[2160] = `CIPHERTEXT_WIDTH'd5598819;
publickey_row[2161] = `CIPHERTEXT_WIDTH'd11950666;
publickey_row[2162] = `CIPHERTEXT_WIDTH'd16626569;
publickey_row[2163] = `CIPHERTEXT_WIDTH'd10607592;
publickey_row[2164] = `CIPHERTEXT_WIDTH'd6209664;
publickey_row[2165] = `CIPHERTEXT_WIDTH'd29631;
publickey_row[2166] = `CIPHERTEXT_WIDTH'd2779165;
publickey_row[2167] = `CIPHERTEXT_WIDTH'd8618377;
publickey_row[2168] = `CIPHERTEXT_WIDTH'd1551559;
publickey_row[2169] = `CIPHERTEXT_WIDTH'd3102603;
publickey_row[2170] = `CIPHERTEXT_WIDTH'd74314;
publickey_row[2171] = `CIPHERTEXT_WIDTH'd5595509;
publickey_row[2172] = `CIPHERTEXT_WIDTH'd16165494;
publickey_row[2173] = `CIPHERTEXT_WIDTH'd8587214;
publickey_row[2174] = `CIPHERTEXT_WIDTH'd9088803;
publickey_row[2175] = `CIPHERTEXT_WIDTH'd1499420;
publickey_row[2176] = `CIPHERTEXT_WIDTH'd10826262;
publickey_row[2177] = `CIPHERTEXT_WIDTH'd15843253;
publickey_row[2178] = `CIPHERTEXT_WIDTH'd9674138;
publickey_row[2179] = `CIPHERTEXT_WIDTH'd8069949;
publickey_row[2180] = `CIPHERTEXT_WIDTH'd15521824;
publickey_row[2181] = `CIPHERTEXT_WIDTH'd14142958;
publickey_row[2182] = `CIPHERTEXT_WIDTH'd13474097;
publickey_row[2183] = `CIPHERTEXT_WIDTH'd6589770;
publickey_row[2184] = `CIPHERTEXT_WIDTH'd14645579;
publickey_row[2185] = `CIPHERTEXT_WIDTH'd7373899;
publickey_row[2186] = `CIPHERTEXT_WIDTH'd15578659;
publickey_row[2187] = `CIPHERTEXT_WIDTH'd5980249;
publickey_row[2188] = `CIPHERTEXT_WIDTH'd14424077;
publickey_row[2189] = `CIPHERTEXT_WIDTH'd8715956;
publickey_row[2190] = `CIPHERTEXT_WIDTH'd10160568;
publickey_row[2191] = `CIPHERTEXT_WIDTH'd1228001;
publickey_row[2192] = `CIPHERTEXT_WIDTH'd5323345;
publickey_row[2193] = `CIPHERTEXT_WIDTH'd7562542;
publickey_row[2194] = `CIPHERTEXT_WIDTH'd15607142;
publickey_row[2195] = `CIPHERTEXT_WIDTH'd12961893;
publickey_row[2196] = `CIPHERTEXT_WIDTH'd12678971;
publickey_row[2197] = `CIPHERTEXT_WIDTH'd4586292;
publickey_row[2198] = `CIPHERTEXT_WIDTH'd15215503;
publickey_row[2199] = `CIPHERTEXT_WIDTH'd6713827;
publickey_row[2200] = `CIPHERTEXT_WIDTH'd11211062;
publickey_row[2201] = `CIPHERTEXT_WIDTH'd4281534;
publickey_row[2202] = `CIPHERTEXT_WIDTH'd1429032;
publickey_row[2203] = `CIPHERTEXT_WIDTH'd12945967;
publickey_row[2204] = `CIPHERTEXT_WIDTH'd6684858;
publickey_row[2205] = `CIPHERTEXT_WIDTH'd10130600;
publickey_row[2206] = `CIPHERTEXT_WIDTH'd10072229;
publickey_row[2207] = `CIPHERTEXT_WIDTH'd12242288;
publickey_row[2208] = `CIPHERTEXT_WIDTH'd10299474;
publickey_row[2209] = `CIPHERTEXT_WIDTH'd8547380;
publickey_row[2210] = `CIPHERTEXT_WIDTH'd10161771;
publickey_row[2211] = `CIPHERTEXT_WIDTH'd11956648;
publickey_row[2212] = `CIPHERTEXT_WIDTH'd4806344;
publickey_row[2213] = `CIPHERTEXT_WIDTH'd8506501;
publickey_row[2214] = `CIPHERTEXT_WIDTH'd5988066;
publickey_row[2215] = `CIPHERTEXT_WIDTH'd8951533;
publickey_row[2216] = `CIPHERTEXT_WIDTH'd15138268;
publickey_row[2217] = `CIPHERTEXT_WIDTH'd4786087;
publickey_row[2218] = `CIPHERTEXT_WIDTH'd12752877;
publickey_row[2219] = `CIPHERTEXT_WIDTH'd5440582;
publickey_row[2220] = `CIPHERTEXT_WIDTH'd11781742;
publickey_row[2221] = `CIPHERTEXT_WIDTH'd6450361;
publickey_row[2222] = `CIPHERTEXT_WIDTH'd16689465;
publickey_row[2223] = `CIPHERTEXT_WIDTH'd12412749;
publickey_row[2224] = `CIPHERTEXT_WIDTH'd16462036;
publickey_row[2225] = `CIPHERTEXT_WIDTH'd8787022;
publickey_row[2226] = `CIPHERTEXT_WIDTH'd15538115;
publickey_row[2227] = `CIPHERTEXT_WIDTH'd200674;
publickey_row[2228] = `CIPHERTEXT_WIDTH'd8374429;
publickey_row[2229] = `CIPHERTEXT_WIDTH'd875792;
publickey_row[2230] = `CIPHERTEXT_WIDTH'd4816717;
publickey_row[2231] = `CIPHERTEXT_WIDTH'd6806600;
publickey_row[2232] = `CIPHERTEXT_WIDTH'd5051780;
publickey_row[2233] = `CIPHERTEXT_WIDTH'd27233;
publickey_row[2234] = `CIPHERTEXT_WIDTH'd14135955;
publickey_row[2235] = `CIPHERTEXT_WIDTH'd15090376;
publickey_row[2236] = `CIPHERTEXT_WIDTH'd4063252;
publickey_row[2237] = `CIPHERTEXT_WIDTH'd12951850;
publickey_row[2238] = `CIPHERTEXT_WIDTH'd3637765;
publickey_row[2239] = `CIPHERTEXT_WIDTH'd11297344;
publickey_row[2240] = `CIPHERTEXT_WIDTH'd10027664;
publickey_row[2241] = `CIPHERTEXT_WIDTH'd8729257;
publickey_row[2242] = `CIPHERTEXT_WIDTH'd14022112;
publickey_row[2243] = `CIPHERTEXT_WIDTH'd3815706;
publickey_row[2244] = `CIPHERTEXT_WIDTH'd4222526;
publickey_row[2245] = `CIPHERTEXT_WIDTH'd14273634;
publickey_row[2246] = `CIPHERTEXT_WIDTH'd1525990;
publickey_row[2247] = `CIPHERTEXT_WIDTH'd3454458;
publickey_row[2248] = `CIPHERTEXT_WIDTH'd3196806;
publickey_row[2249] = `CIPHERTEXT_WIDTH'd2098038;
publickey_row[2250] = `CIPHERTEXT_WIDTH'd14444258;
publickey_row[2251] = `CIPHERTEXT_WIDTH'd8990561;
publickey_row[2252] = `CIPHERTEXT_WIDTH'd2061446;
publickey_row[2253] = `CIPHERTEXT_WIDTH'd7786532;
publickey_row[2254] = `CIPHERTEXT_WIDTH'd10067220;
publickey_row[2255] = `CIPHERTEXT_WIDTH'd16223879;
publickey_row[2256] = `CIPHERTEXT_WIDTH'd4439271;
publickey_row[2257] = `CIPHERTEXT_WIDTH'd13241737;
publickey_row[2258] = `CIPHERTEXT_WIDTH'd9055497;
publickey_row[2259] = `CIPHERTEXT_WIDTH'd10158896;
publickey_row[2260] = `CIPHERTEXT_WIDTH'd8613564;
publickey_row[2261] = `CIPHERTEXT_WIDTH'd11915208;
publickey_row[2262] = `CIPHERTEXT_WIDTH'd1744811;
publickey_row[2263] = `CIPHERTEXT_WIDTH'd7152334;
publickey_row[2264] = `CIPHERTEXT_WIDTH'd8095794;
publickey_row[2265] = `CIPHERTEXT_WIDTH'd13226736;
publickey_row[2266] = `CIPHERTEXT_WIDTH'd13984805;
publickey_row[2267] = `CIPHERTEXT_WIDTH'd14566242;
publickey_row[2268] = `CIPHERTEXT_WIDTH'd14956638;
publickey_row[2269] = `CIPHERTEXT_WIDTH'd5004196;
publickey_row[2270] = `CIPHERTEXT_WIDTH'd7504894;
publickey_row[2271] = `CIPHERTEXT_WIDTH'd4382397;
publickey_row[2272] = `CIPHERTEXT_WIDTH'd2674291;
publickey_row[2273] = `CIPHERTEXT_WIDTH'd9436289;
publickey_row[2274] = `CIPHERTEXT_WIDTH'd12142;
publickey_row[2275] = `CIPHERTEXT_WIDTH'd7835431;
publickey_row[2276] = `CIPHERTEXT_WIDTH'd9017485;
publickey_row[2277] = `CIPHERTEXT_WIDTH'd1566790;
publickey_row[2278] = `CIPHERTEXT_WIDTH'd5392971;
publickey_row[2279] = `CIPHERTEXT_WIDTH'd12313030;
publickey_row[2280] = `CIPHERTEXT_WIDTH'd11433934;
publickey_row[2281] = `CIPHERTEXT_WIDTH'd3339345;
publickey_row[2282] = `CIPHERTEXT_WIDTH'd10993389;
publickey_row[2283] = `CIPHERTEXT_WIDTH'd5855873;
publickey_row[2284] = `CIPHERTEXT_WIDTH'd1141550;
publickey_row[2285] = `CIPHERTEXT_WIDTH'd509089;
publickey_row[2286] = `CIPHERTEXT_WIDTH'd3459212;
publickey_row[2287] = `CIPHERTEXT_WIDTH'd13114141;
publickey_row[2288] = `CIPHERTEXT_WIDTH'd9989281;
publickey_row[2289] = `CIPHERTEXT_WIDTH'd5802235;
publickey_row[2290] = `CIPHERTEXT_WIDTH'd5282952;
publickey_row[2291] = `CIPHERTEXT_WIDTH'd13900333;
publickey_row[2292] = `CIPHERTEXT_WIDTH'd4537918;
publickey_row[2293] = `CIPHERTEXT_WIDTH'd1636596;
publickey_row[2294] = `CIPHERTEXT_WIDTH'd14969688;
publickey_row[2295] = `CIPHERTEXT_WIDTH'd9811890;
publickey_row[2296] = `CIPHERTEXT_WIDTH'd13935618;
publickey_row[2297] = `CIPHERTEXT_WIDTH'd4707094;
publickey_row[2298] = `CIPHERTEXT_WIDTH'd9708726;
publickey_row[2299] = `CIPHERTEXT_WIDTH'd685557;
publickey_row[2300] = `CIPHERTEXT_WIDTH'd2887038;
publickey_row[2301] = `CIPHERTEXT_WIDTH'd14139607;
publickey_row[2302] = `CIPHERTEXT_WIDTH'd10159212;
publickey_row[2303] = `CIPHERTEXT_WIDTH'd7382021;
publickey_row[2304] = `CIPHERTEXT_WIDTH'd8271807;
publickey_row[2305] = `CIPHERTEXT_WIDTH'd714477;
publickey_row[2306] = `CIPHERTEXT_WIDTH'd15727516;
publickey_row[2307] = `CIPHERTEXT_WIDTH'd15339558;
publickey_row[2308] = `CIPHERTEXT_WIDTH'd4658428;
publickey_row[2309] = `CIPHERTEXT_WIDTH'd8073803;
publickey_row[2310] = `CIPHERTEXT_WIDTH'd4417391;
publickey_row[2311] = `CIPHERTEXT_WIDTH'd8899085;
publickey_row[2312] = `CIPHERTEXT_WIDTH'd1937286;
publickey_row[2313] = `CIPHERTEXT_WIDTH'd3279265;
publickey_row[2314] = `CIPHERTEXT_WIDTH'd10562522;
publickey_row[2315] = `CIPHERTEXT_WIDTH'd497390;
publickey_row[2316] = `CIPHERTEXT_WIDTH'd15662318;
publickey_row[2317] = `CIPHERTEXT_WIDTH'd16644432;
publickey_row[2318] = `CIPHERTEXT_WIDTH'd1452176;
publickey_row[2319] = `CIPHERTEXT_WIDTH'd1578423;
publickey_row[2320] = `CIPHERTEXT_WIDTH'd11841228;
publickey_row[2321] = `CIPHERTEXT_WIDTH'd685102;
publickey_row[2322] = `CIPHERTEXT_WIDTH'd12240055;
publickey_row[2323] = `CIPHERTEXT_WIDTH'd3896249;
publickey_row[2324] = `CIPHERTEXT_WIDTH'd4901657;
publickey_row[2325] = `CIPHERTEXT_WIDTH'd2987144;
publickey_row[2326] = `CIPHERTEXT_WIDTH'd16439399;
publickey_row[2327] = `CIPHERTEXT_WIDTH'd8294903;
publickey_row[2328] = `CIPHERTEXT_WIDTH'd10378654;
publickey_row[2329] = `CIPHERTEXT_WIDTH'd12378365;
publickey_row[2330] = `CIPHERTEXT_WIDTH'd5274358;
publickey_row[2331] = `CIPHERTEXT_WIDTH'd9324526;
publickey_row[2332] = `CIPHERTEXT_WIDTH'd1493122;
publickey_row[2333] = `CIPHERTEXT_WIDTH'd8447736;
publickey_row[2334] = `CIPHERTEXT_WIDTH'd56565;
publickey_row[2335] = `CIPHERTEXT_WIDTH'd7296336;
publickey_row[2336] = `CIPHERTEXT_WIDTH'd8672039;
publickey_row[2337] = `CIPHERTEXT_WIDTH'd4220670;
publickey_row[2338] = `CIPHERTEXT_WIDTH'd16654192;
publickey_row[2339] = `CIPHERTEXT_WIDTH'd7680461;
publickey_row[2340] = `CIPHERTEXT_WIDTH'd8597699;
publickey_row[2341] = `CIPHERTEXT_WIDTH'd1874364;
publickey_row[2342] = `CIPHERTEXT_WIDTH'd10289025;
publickey_row[2343] = `CIPHERTEXT_WIDTH'd6982717;
publickey_row[2344] = `CIPHERTEXT_WIDTH'd6016823;
publickey_row[2345] = `CIPHERTEXT_WIDTH'd10533160;
publickey_row[2346] = `CIPHERTEXT_WIDTH'd5227634;
publickey_row[2347] = `CIPHERTEXT_WIDTH'd3210370;
publickey_row[2348] = `CIPHERTEXT_WIDTH'd12376382;
publickey_row[2349] = `CIPHERTEXT_WIDTH'd7515753;
publickey_row[2350] = `CIPHERTEXT_WIDTH'd16133760;
publickey_row[2351] = `CIPHERTEXT_WIDTH'd4893445;
publickey_row[2352] = `CIPHERTEXT_WIDTH'd8654330;
publickey_row[2353] = `CIPHERTEXT_WIDTH'd7117123;
publickey_row[2354] = `CIPHERTEXT_WIDTH'd1779597;
publickey_row[2355] = `CIPHERTEXT_WIDTH'd1499046;
publickey_row[2356] = `CIPHERTEXT_WIDTH'd12229185;
publickey_row[2357] = `CIPHERTEXT_WIDTH'd6546407;
publickey_row[2358] = `CIPHERTEXT_WIDTH'd8276210;
publickey_row[2359] = `CIPHERTEXT_WIDTH'd8259099;
publickey_row[2360] = `CIPHERTEXT_WIDTH'd11944392;
publickey_row[2361] = `CIPHERTEXT_WIDTH'd12989532;
publickey_row[2362] = `CIPHERTEXT_WIDTH'd4777891;
publickey_row[2363] = `CIPHERTEXT_WIDTH'd5145383;
publickey_row[2364] = `CIPHERTEXT_WIDTH'd12752651;
publickey_row[2365] = `CIPHERTEXT_WIDTH'd2172243;
publickey_row[2366] = `CIPHERTEXT_WIDTH'd15229530;
publickey_row[2367] = `CIPHERTEXT_WIDTH'd13941077;
publickey_row[2368] = `CIPHERTEXT_WIDTH'd6660711;
publickey_row[2369] = `CIPHERTEXT_WIDTH'd12872510;
publickey_row[2370] = `CIPHERTEXT_WIDTH'd9907964;
publickey_row[2371] = `CIPHERTEXT_WIDTH'd16743409;
publickey_row[2372] = `CIPHERTEXT_WIDTH'd2322788;
publickey_row[2373] = `CIPHERTEXT_WIDTH'd184821;
publickey_row[2374] = `CIPHERTEXT_WIDTH'd5429194;
publickey_row[2375] = `CIPHERTEXT_WIDTH'd13500313;
publickey_row[2376] = `CIPHERTEXT_WIDTH'd8476461;
publickey_row[2377] = `CIPHERTEXT_WIDTH'd9548227;
publickey_row[2378] = `CIPHERTEXT_WIDTH'd15705509;
publickey_row[2379] = `CIPHERTEXT_WIDTH'd6569703;
publickey_row[2380] = `CIPHERTEXT_WIDTH'd201860;
publickey_row[2381] = `CIPHERTEXT_WIDTH'd4341716;
publickey_row[2382] = `CIPHERTEXT_WIDTH'd10991356;
publickey_row[2383] = `CIPHERTEXT_WIDTH'd6714114;
publickey_row[2384] = `CIPHERTEXT_WIDTH'd2746323;
publickey_row[2385] = `CIPHERTEXT_WIDTH'd16556153;
publickey_row[2386] = `CIPHERTEXT_WIDTH'd1792900;
publickey_row[2387] = `CIPHERTEXT_WIDTH'd6036655;
publickey_row[2388] = `CIPHERTEXT_WIDTH'd9677147;
publickey_row[2389] = `CIPHERTEXT_WIDTH'd3275907;
publickey_row[2390] = `CIPHERTEXT_WIDTH'd12045199;
publickey_row[2391] = `CIPHERTEXT_WIDTH'd16621955;
publickey_row[2392] = `CIPHERTEXT_WIDTH'd6073110;
publickey_row[2393] = `CIPHERTEXT_WIDTH'd4079131;
publickey_row[2394] = `CIPHERTEXT_WIDTH'd5762735;
publickey_row[2395] = `CIPHERTEXT_WIDTH'd15601779;
publickey_row[2396] = `CIPHERTEXT_WIDTH'd3253645;
publickey_row[2397] = `CIPHERTEXT_WIDTH'd5274248;
publickey_row[2398] = `CIPHERTEXT_WIDTH'd7556194;
publickey_row[2399] = `CIPHERTEXT_WIDTH'd1358154;
publickey_row[2400] = `CIPHERTEXT_WIDTH'd4640019;
publickey_row[2401] = `CIPHERTEXT_WIDTH'd9859711;
publickey_row[2402] = `CIPHERTEXT_WIDTH'd15654640;
publickey_row[2403] = `CIPHERTEXT_WIDTH'd6396420;
publickey_row[2404] = `CIPHERTEXT_WIDTH'd9609553;
publickey_row[2405] = `CIPHERTEXT_WIDTH'd7469487;
publickey_row[2406] = `CIPHERTEXT_WIDTH'd9751935;
publickey_row[2407] = `CIPHERTEXT_WIDTH'd14659735;
publickey_row[2408] = `CIPHERTEXT_WIDTH'd15472189;
publickey_row[2409] = `CIPHERTEXT_WIDTH'd4122508;
publickey_row[2410] = `CIPHERTEXT_WIDTH'd11175787;
publickey_row[2411] = `CIPHERTEXT_WIDTH'd16399957;
publickey_row[2412] = `CIPHERTEXT_WIDTH'd13172164;
publickey_row[2413] = `CIPHERTEXT_WIDTH'd14911067;
publickey_row[2414] = `CIPHERTEXT_WIDTH'd9676411;
publickey_row[2415] = `CIPHERTEXT_WIDTH'd16741079;
publickey_row[2416] = `CIPHERTEXT_WIDTH'd14003176;
publickey_row[2417] = `CIPHERTEXT_WIDTH'd15656863;
publickey_row[2418] = `CIPHERTEXT_WIDTH'd14527980;
publickey_row[2419] = `CIPHERTEXT_WIDTH'd8249437;
publickey_row[2420] = `CIPHERTEXT_WIDTH'd10681408;
publickey_row[2421] = `CIPHERTEXT_WIDTH'd936612;
publickey_row[2422] = `CIPHERTEXT_WIDTH'd828098;
publickey_row[2423] = `CIPHERTEXT_WIDTH'd484748;
publickey_row[2424] = `CIPHERTEXT_WIDTH'd13309870;
publickey_row[2425] = `CIPHERTEXT_WIDTH'd363431;
publickey_row[2426] = `CIPHERTEXT_WIDTH'd14615958;
publickey_row[2427] = `CIPHERTEXT_WIDTH'd15484964;
publickey_row[2428] = `CIPHERTEXT_WIDTH'd3495075;
publickey_row[2429] = `CIPHERTEXT_WIDTH'd5700510;
publickey_row[2430] = `CIPHERTEXT_WIDTH'd9173849;
publickey_row[2431] = `CIPHERTEXT_WIDTH'd13333921;
publickey_row[2432] = `CIPHERTEXT_WIDTH'd15185528;
publickey_row[2433] = `CIPHERTEXT_WIDTH'd12191111;
publickey_row[2434] = `CIPHERTEXT_WIDTH'd15535922;
publickey_row[2435] = `CIPHERTEXT_WIDTH'd4949579;
publickey_row[2436] = `CIPHERTEXT_WIDTH'd10182404;
publickey_row[2437] = `CIPHERTEXT_WIDTH'd14957653;
publickey_row[2438] = `CIPHERTEXT_WIDTH'd8427878;
publickey_row[2439] = `CIPHERTEXT_WIDTH'd3686855;
publickey_row[2440] = `CIPHERTEXT_WIDTH'd1702073;
publickey_row[2441] = `CIPHERTEXT_WIDTH'd820390;
publickey_row[2442] = `CIPHERTEXT_WIDTH'd16305505;
publickey_row[2443] = `CIPHERTEXT_WIDTH'd8607179;
publickey_row[2444] = `CIPHERTEXT_WIDTH'd10474055;
publickey_row[2445] = `CIPHERTEXT_WIDTH'd5502669;
publickey_row[2446] = `CIPHERTEXT_WIDTH'd1774529;
publickey_row[2447] = `CIPHERTEXT_WIDTH'd4562182;
publickey_row[2448] = `CIPHERTEXT_WIDTH'd2386564;
publickey_row[2449] = `CIPHERTEXT_WIDTH'd1150179;
publickey_row[2450] = `CIPHERTEXT_WIDTH'd13930613;
publickey_row[2451] = `CIPHERTEXT_WIDTH'd15470266;
publickey_row[2452] = `CIPHERTEXT_WIDTH'd13221123;
publickey_row[2453] = `CIPHERTEXT_WIDTH'd14396186;
publickey_row[2454] = `CIPHERTEXT_WIDTH'd10826784;
publickey_row[2455] = `CIPHERTEXT_WIDTH'd9921860;
publickey_row[2456] = `CIPHERTEXT_WIDTH'd4378735;
publickey_row[2457] = `CIPHERTEXT_WIDTH'd3026167;
publickey_row[2458] = `CIPHERTEXT_WIDTH'd14900698;
publickey_row[2459] = `CIPHERTEXT_WIDTH'd15368961;
publickey_row[2460] = `CIPHERTEXT_WIDTH'd9208132;
publickey_row[2461] = `CIPHERTEXT_WIDTH'd15262115;
publickey_row[2462] = `CIPHERTEXT_WIDTH'd14913710;
publickey_row[2463] = `CIPHERTEXT_WIDTH'd4128337;
publickey_row[2464] = `CIPHERTEXT_WIDTH'd16720089;
publickey_row[2465] = `CIPHERTEXT_WIDTH'd7312759;
publickey_row[2466] = `CIPHERTEXT_WIDTH'd12324945;
publickey_row[2467] = `CIPHERTEXT_WIDTH'd1492186;
publickey_row[2468] = `CIPHERTEXT_WIDTH'd6442079;
publickey_row[2469] = `CIPHERTEXT_WIDTH'd13708046;
publickey_row[2470] = `CIPHERTEXT_WIDTH'd14750882;
publickey_row[2471] = `CIPHERTEXT_WIDTH'd6907996;
publickey_row[2472] = `CIPHERTEXT_WIDTH'd7473732;
publickey_row[2473] = `CIPHERTEXT_WIDTH'd6927912;
publickey_row[2474] = `CIPHERTEXT_WIDTH'd751958;
publickey_row[2475] = `CIPHERTEXT_WIDTH'd12094611;
publickey_row[2476] = `CIPHERTEXT_WIDTH'd16769866;
publickey_row[2477] = `CIPHERTEXT_WIDTH'd15429407;
publickey_row[2478] = `CIPHERTEXT_WIDTH'd1742970;
publickey_row[2479] = `CIPHERTEXT_WIDTH'd14737909;
publickey_row[2480] = `CIPHERTEXT_WIDTH'd15616790;
publickey_row[2481] = `CIPHERTEXT_WIDTH'd1866683;
publickey_row[2482] = `CIPHERTEXT_WIDTH'd10061224;
publickey_row[2483] = `CIPHERTEXT_WIDTH'd15709943;
publickey_row[2484] = `CIPHERTEXT_WIDTH'd7553813;
publickey_row[2485] = `CIPHERTEXT_WIDTH'd1479333;
publickey_row[2486] = `CIPHERTEXT_WIDTH'd13647342;
publickey_row[2487] = `CIPHERTEXT_WIDTH'd4587261;
publickey_row[2488] = `CIPHERTEXT_WIDTH'd8759734;
publickey_row[2489] = `CIPHERTEXT_WIDTH'd1201014;
publickey_row[2490] = `CIPHERTEXT_WIDTH'd6945265;
publickey_row[2491] = `CIPHERTEXT_WIDTH'd9240004;
publickey_row[2492] = `CIPHERTEXT_WIDTH'd10280518;
publickey_row[2493] = `CIPHERTEXT_WIDTH'd2383377;
publickey_row[2494] = `CIPHERTEXT_WIDTH'd10164475;
publickey_row[2495] = `CIPHERTEXT_WIDTH'd3858648;
publickey_row[2496] = `CIPHERTEXT_WIDTH'd12663236;
publickey_row[2497] = `CIPHERTEXT_WIDTH'd13914259;
publickey_row[2498] = `CIPHERTEXT_WIDTH'd4057328;
publickey_row[2499] = `CIPHERTEXT_WIDTH'd12208871;
publickey_row[2500] = `CIPHERTEXT_WIDTH'd5530527;
publickey_row[2501] = `CIPHERTEXT_WIDTH'd6655280;
publickey_row[2502] = `CIPHERTEXT_WIDTH'd4789541;
publickey_row[2503] = `CIPHERTEXT_WIDTH'd11973585;
publickey_row[2504] = `CIPHERTEXT_WIDTH'd3998714;
publickey_row[2505] = `CIPHERTEXT_WIDTH'd15340438;
publickey_row[2506] = `CIPHERTEXT_WIDTH'd4894778;
publickey_row[2507] = `CIPHERTEXT_WIDTH'd2479337;
publickey_row[2508] = `CIPHERTEXT_WIDTH'd13572069;
publickey_row[2509] = `CIPHERTEXT_WIDTH'd6644977;
publickey_row[2510] = `CIPHERTEXT_WIDTH'd14049420;
publickey_row[2511] = `CIPHERTEXT_WIDTH'd12237628;
publickey_row[2512] = `CIPHERTEXT_WIDTH'd13020520;
publickey_row[2513] = `CIPHERTEXT_WIDTH'd10562062;
publickey_row[2514] = `CIPHERTEXT_WIDTH'd14131323;
publickey_row[2515] = `CIPHERTEXT_WIDTH'd8729614;
publickey_row[2516] = `CIPHERTEXT_WIDTH'd12543946;
publickey_row[2517] = `CIPHERTEXT_WIDTH'd14671417;
publickey_row[2518] = `CIPHERTEXT_WIDTH'd3262908;
publickey_row[2519] = `CIPHERTEXT_WIDTH'd2585620;
publickey_row[2520] = `CIPHERTEXT_WIDTH'd10529653;
publickey_row[2521] = `CIPHERTEXT_WIDTH'd14777593;
publickey_row[2522] = `CIPHERTEXT_WIDTH'd5578958;
publickey_row[2523] = `CIPHERTEXT_WIDTH'd1843167;
publickey_row[2524] = `CIPHERTEXT_WIDTH'd9700158;
publickey_row[2525] = `CIPHERTEXT_WIDTH'd12671865;
publickey_row[2526] = `CIPHERTEXT_WIDTH'd963231;
publickey_row[2527] = `CIPHERTEXT_WIDTH'd4001173;
publickey_row[2528] = `CIPHERTEXT_WIDTH'd2690008;
publickey_row[2529] = `CIPHERTEXT_WIDTH'd5860138;
publickey_row[2530] = `CIPHERTEXT_WIDTH'd12677126;
publickey_row[2531] = `CIPHERTEXT_WIDTH'd876174;
publickey_row[2532] = `CIPHERTEXT_WIDTH'd5794704;
publickey_row[2533] = `CIPHERTEXT_WIDTH'd10273804;
publickey_row[2534] = `CIPHERTEXT_WIDTH'd3555482;
publickey_row[2535] = `CIPHERTEXT_WIDTH'd6261838;
publickey_row[2536] = `CIPHERTEXT_WIDTH'd3566251;
publickey_row[2537] = `CIPHERTEXT_WIDTH'd1352324;
publickey_row[2538] = `CIPHERTEXT_WIDTH'd148982;
publickey_row[2539] = `CIPHERTEXT_WIDTH'd2353229;
publickey_row[2540] = `CIPHERTEXT_WIDTH'd9367958;
publickey_row[2541] = `CIPHERTEXT_WIDTH'd15748190;
publickey_row[2542] = `CIPHERTEXT_WIDTH'd8312687;
publickey_row[2543] = `CIPHERTEXT_WIDTH'd8076765;
publickey_row[2544] = `CIPHERTEXT_WIDTH'd12870084;
publickey_row[2545] = `CIPHERTEXT_WIDTH'd8953525;
publickey_row[2546] = `CIPHERTEXT_WIDTH'd11495621;
publickey_row[2547] = `CIPHERTEXT_WIDTH'd3390322;
publickey_row[2548] = `CIPHERTEXT_WIDTH'd16527861;
publickey_row[2549] = `CIPHERTEXT_WIDTH'd515754;
publickey_row[2550] = `CIPHERTEXT_WIDTH'd5983102;
publickey_row[2551] = `CIPHERTEXT_WIDTH'd14003881;
publickey_row[2552] = `CIPHERTEXT_WIDTH'd15256338;
publickey_row[2553] = `CIPHERTEXT_WIDTH'd3621016;
publickey_row[2554] = `CIPHERTEXT_WIDTH'd9181706;
publickey_row[2555] = `CIPHERTEXT_WIDTH'd4841803;
publickey_row[2556] = `CIPHERTEXT_WIDTH'd14912881;
publickey_row[2557] = `CIPHERTEXT_WIDTH'd8412655;
publickey_row[2558] = `CIPHERTEXT_WIDTH'd12482349;
publickey_row[2559] = `CIPHERTEXT_WIDTH'd16158095;
publickey_row[2560] = `CIPHERTEXT_WIDTH'd7150802;
publickey_row[2561] = `CIPHERTEXT_WIDTH'd9090408;
publickey_row[2562] = `CIPHERTEXT_WIDTH'd5845540;
publickey_row[2563] = `CIPHERTEXT_WIDTH'd7033591;
publickey_row[2564] = `CIPHERTEXT_WIDTH'd3195610;
publickey_row[2565] = `CIPHERTEXT_WIDTH'd12637747;
publickey_row[2566] = `CIPHERTEXT_WIDTH'd6538229;
publickey_row[2567] = `CIPHERTEXT_WIDTH'd1154760;
publickey_row[2568] = `CIPHERTEXT_WIDTH'd11350817;
publickey_row[2569] = `CIPHERTEXT_WIDTH'd1342269;
publickey_row[2570] = `CIPHERTEXT_WIDTH'd10713558;
publickey_row[2571] = `CIPHERTEXT_WIDTH'd16656135;
publickey_row[2572] = `CIPHERTEXT_WIDTH'd960424;
publickey_row[2573] = `CIPHERTEXT_WIDTH'd2088742;
publickey_row[2574] = `CIPHERTEXT_WIDTH'd15830086;
publickey_row[2575] = `CIPHERTEXT_WIDTH'd12965096;
publickey_row[2576] = `CIPHERTEXT_WIDTH'd3481884;
publickey_row[2577] = `CIPHERTEXT_WIDTH'd10644233;
publickey_row[2578] = `CIPHERTEXT_WIDTH'd4324164;
publickey_row[2579] = `CIPHERTEXT_WIDTH'd1280678;
publickey_row[2580] = `CIPHERTEXT_WIDTH'd13499983;
publickey_row[2581] = `CIPHERTEXT_WIDTH'd14071856;
publickey_row[2582] = `CIPHERTEXT_WIDTH'd5058142;
publickey_row[2583] = `CIPHERTEXT_WIDTH'd7661349;
publickey_row[2584] = `CIPHERTEXT_WIDTH'd4312213;
publickey_row[2585] = `CIPHERTEXT_WIDTH'd2116300;
publickey_row[2586] = `CIPHERTEXT_WIDTH'd7020308;
publickey_row[2587] = `CIPHERTEXT_WIDTH'd11359604;
publickey_row[2588] = `CIPHERTEXT_WIDTH'd9414702;
publickey_row[2589] = `CIPHERTEXT_WIDTH'd13450223;
publickey_row[2590] = `CIPHERTEXT_WIDTH'd3839961;
publickey_row[2591] = `CIPHERTEXT_WIDTH'd4244972;
publickey_row[2592] = `CIPHERTEXT_WIDTH'd1934743;
publickey_row[2593] = `CIPHERTEXT_WIDTH'd16322981;
publickey_row[2594] = `CIPHERTEXT_WIDTH'd3115682;
publickey_row[2595] = `CIPHERTEXT_WIDTH'd12032923;
publickey_row[2596] = `CIPHERTEXT_WIDTH'd1766167;
publickey_row[2597] = `CIPHERTEXT_WIDTH'd12032704;
publickey_row[2598] = `CIPHERTEXT_WIDTH'd11178940;
publickey_row[2599] = `CIPHERTEXT_WIDTH'd8928809;
publickey_row[2600] = `CIPHERTEXT_WIDTH'd4225997;
publickey_row[2601] = `CIPHERTEXT_WIDTH'd858587;
publickey_row[2602] = `CIPHERTEXT_WIDTH'd444724;
publickey_row[2603] = `CIPHERTEXT_WIDTH'd15752369;
publickey_row[2604] = `CIPHERTEXT_WIDTH'd1539395;
publickey_row[2605] = `CIPHERTEXT_WIDTH'd938862;
publickey_row[2606] = `CIPHERTEXT_WIDTH'd8005519;
publickey_row[2607] = `CIPHERTEXT_WIDTH'd8872278;
publickey_row[2608] = `CIPHERTEXT_WIDTH'd5461580;
publickey_row[2609] = `CIPHERTEXT_WIDTH'd7656573;
publickey_row[2610] = `CIPHERTEXT_WIDTH'd4007226;
publickey_row[2611] = `CIPHERTEXT_WIDTH'd13119420;
publickey_row[2612] = `CIPHERTEXT_WIDTH'd5676138;
publickey_row[2613] = `CIPHERTEXT_WIDTH'd16424367;
publickey_row[2614] = `CIPHERTEXT_WIDTH'd16316001;
publickey_row[2615] = `CIPHERTEXT_WIDTH'd13999530;
publickey_row[2616] = `CIPHERTEXT_WIDTH'd7586509;
publickey_row[2617] = `CIPHERTEXT_WIDTH'd9469;
publickey_row[2618] = `CIPHERTEXT_WIDTH'd14012443;
publickey_row[2619] = `CIPHERTEXT_WIDTH'd7354018;
publickey_row[2620] = `CIPHERTEXT_WIDTH'd1141673;
publickey_row[2621] = `CIPHERTEXT_WIDTH'd7572232;
publickey_row[2622] = `CIPHERTEXT_WIDTH'd14891716;
publickey_row[2623] = `CIPHERTEXT_WIDTH'd10757105;
publickey_row[2624] = `CIPHERTEXT_WIDTH'd14770802;
publickey_row[2625] = `CIPHERTEXT_WIDTH'd3436187;
publickey_row[2626] = `CIPHERTEXT_WIDTH'd14078423;
publickey_row[2627] = `CIPHERTEXT_WIDTH'd2995858;
publickey_row[2628] = `CIPHERTEXT_WIDTH'd9810366;
publickey_row[2629] = `CIPHERTEXT_WIDTH'd13897858;
publickey_row[2630] = `CIPHERTEXT_WIDTH'd1442059;
publickey_row[2631] = `CIPHERTEXT_WIDTH'd3881988;
publickey_row[2632] = `CIPHERTEXT_WIDTH'd4141197;
publickey_row[2633] = `CIPHERTEXT_WIDTH'd8349000;
publickey_row[2634] = `CIPHERTEXT_WIDTH'd12061612;
publickey_row[2635] = `CIPHERTEXT_WIDTH'd582224;
publickey_row[2636] = `CIPHERTEXT_WIDTH'd8102453;
publickey_row[2637] = `CIPHERTEXT_WIDTH'd14325330;
publickey_row[2638] = `CIPHERTEXT_WIDTH'd11353852;
publickey_row[2639] = `CIPHERTEXT_WIDTH'd4170433;
publickey_row[2640] = `CIPHERTEXT_WIDTH'd3051745;
publickey_row[2641] = `CIPHERTEXT_WIDTH'd10144376;
publickey_row[2642] = `CIPHERTEXT_WIDTH'd9886768;
publickey_row[2643] = `CIPHERTEXT_WIDTH'd11727398;
publickey_row[2644] = `CIPHERTEXT_WIDTH'd15865529;
publickey_row[2645] = `CIPHERTEXT_WIDTH'd3761012;
publickey_row[2646] = `CIPHERTEXT_WIDTH'd15666324;
publickey_row[2647] = `CIPHERTEXT_WIDTH'd8261684;
publickey_row[2648] = `CIPHERTEXT_WIDTH'd14469764;
publickey_row[2649] = `CIPHERTEXT_WIDTH'd12361869;
publickey_row[2650] = `CIPHERTEXT_WIDTH'd8781427;
publickey_row[2651] = `CIPHERTEXT_WIDTH'd4501053;
publickey_row[2652] = `CIPHERTEXT_WIDTH'd1674114;
publickey_row[2653] = `CIPHERTEXT_WIDTH'd2756252;
publickey_row[2654] = `CIPHERTEXT_WIDTH'd13562991;
publickey_row[2655] = `CIPHERTEXT_WIDTH'd4383163;
publickey_row[2656] = `CIPHERTEXT_WIDTH'd11471174;
publickey_row[2657] = `CIPHERTEXT_WIDTH'd15921426;
publickey_row[2658] = `CIPHERTEXT_WIDTH'd8789936;
publickey_row[2659] = `CIPHERTEXT_WIDTH'd10006795;
publickey_row[2660] = `CIPHERTEXT_WIDTH'd2487935;
publickey_row[2661] = `CIPHERTEXT_WIDTH'd12448210;
publickey_row[2662] = `CIPHERTEXT_WIDTH'd13687360;
publickey_row[2663] = `CIPHERTEXT_WIDTH'd7802069;
publickey_row[2664] = `CIPHERTEXT_WIDTH'd1550647;
publickey_row[2665] = `CIPHERTEXT_WIDTH'd2680643;
publickey_row[2666] = `CIPHERTEXT_WIDTH'd912536;
publickey_row[2667] = `CIPHERTEXT_WIDTH'd11719611;
publickey_row[2668] = `CIPHERTEXT_WIDTH'd16751651;
publickey_row[2669] = `CIPHERTEXT_WIDTH'd16383822;
publickey_row[2670] = `CIPHERTEXT_WIDTH'd11234887;
publickey_row[2671] = `CIPHERTEXT_WIDTH'd12282154;
publickey_row[2672] = `CIPHERTEXT_WIDTH'd15485132;
publickey_row[2673] = `CIPHERTEXT_WIDTH'd12362174;
publickey_row[2674] = `CIPHERTEXT_WIDTH'd10731762;
publickey_row[2675] = `CIPHERTEXT_WIDTH'd253019;
publickey_row[2676] = `CIPHERTEXT_WIDTH'd11594914;
publickey_row[2677] = `CIPHERTEXT_WIDTH'd12722465;
publickey_row[2678] = `CIPHERTEXT_WIDTH'd441128;
publickey_row[2679] = `CIPHERTEXT_WIDTH'd13036342;
publickey_row[2680] = `CIPHERTEXT_WIDTH'd8211051;
publickey_row[2681] = `CIPHERTEXT_WIDTH'd1110530;
publickey_row[2682] = `CIPHERTEXT_WIDTH'd16399775;
publickey_row[2683] = `CIPHERTEXT_WIDTH'd10725275;
publickey_row[2684] = `CIPHERTEXT_WIDTH'd14409161;
publickey_row[2685] = `CIPHERTEXT_WIDTH'd398457;
publickey_row[2686] = `CIPHERTEXT_WIDTH'd6912439;
publickey_row[2687] = `CIPHERTEXT_WIDTH'd12079626;
publickey_row[2688] = `CIPHERTEXT_WIDTH'd13373481;
publickey_row[2689] = `CIPHERTEXT_WIDTH'd13433330;
publickey_row[2690] = `CIPHERTEXT_WIDTH'd3131757;
publickey_row[2691] = `CIPHERTEXT_WIDTH'd10383950;
publickey_row[2692] = `CIPHERTEXT_WIDTH'd4377595;
publickey_row[2693] = `CIPHERTEXT_WIDTH'd16377329;
publickey_row[2694] = `CIPHERTEXT_WIDTH'd11129370;
publickey_row[2695] = `CIPHERTEXT_WIDTH'd4847400;
publickey_row[2696] = `CIPHERTEXT_WIDTH'd1986525;
publickey_row[2697] = `CIPHERTEXT_WIDTH'd888024;
publickey_row[2698] = `CIPHERTEXT_WIDTH'd4935188;
publickey_row[2699] = `CIPHERTEXT_WIDTH'd2960781;
publickey_row[2700] = `CIPHERTEXT_WIDTH'd15092684;
publickey_row[2701] = `CIPHERTEXT_WIDTH'd10262166;
publickey_row[2702] = `CIPHERTEXT_WIDTH'd1201293;
publickey_row[2703] = `CIPHERTEXT_WIDTH'd13861489;
publickey_row[2704] = `CIPHERTEXT_WIDTH'd8376721;
publickey_row[2705] = `CIPHERTEXT_WIDTH'd11818933;
publickey_row[2706] = `CIPHERTEXT_WIDTH'd242770;
publickey_row[2707] = `CIPHERTEXT_WIDTH'd13743947;
publickey_row[2708] = `CIPHERTEXT_WIDTH'd13113004;
publickey_row[2709] = `CIPHERTEXT_WIDTH'd3327497;
publickey_row[2710] = `CIPHERTEXT_WIDTH'd14132213;
publickey_row[2711] = `CIPHERTEXT_WIDTH'd3581310;
publickey_row[2712] = `CIPHERTEXT_WIDTH'd11775943;
publickey_row[2713] = `CIPHERTEXT_WIDTH'd12094305;
publickey_row[2714] = `CIPHERTEXT_WIDTH'd16757010;
publickey_row[2715] = `CIPHERTEXT_WIDTH'd11753213;
publickey_row[2716] = `CIPHERTEXT_WIDTH'd995281;
publickey_row[2717] = `CIPHERTEXT_WIDTH'd15814333;
publickey_row[2718] = `CIPHERTEXT_WIDTH'd5674831;
publickey_row[2719] = `CIPHERTEXT_WIDTH'd1876229;
publickey_row[2720] = `CIPHERTEXT_WIDTH'd8792674;
publickey_row[2721] = `CIPHERTEXT_WIDTH'd2549612;
publickey_row[2722] = `CIPHERTEXT_WIDTH'd13314105;
publickey_row[2723] = `CIPHERTEXT_WIDTH'd14182582;
publickey_row[2724] = `CIPHERTEXT_WIDTH'd13170032;
publickey_row[2725] = `CIPHERTEXT_WIDTH'd13952716;
publickey_row[2726] = `CIPHERTEXT_WIDTH'd4327989;
publickey_row[2727] = `CIPHERTEXT_WIDTH'd10437380;
publickey_row[2728] = `CIPHERTEXT_WIDTH'd7871137;
publickey_row[2729] = `CIPHERTEXT_WIDTH'd3609770;
publickey_row[2730] = `CIPHERTEXT_WIDTH'd11540656;
publickey_row[2731] = `CIPHERTEXT_WIDTH'd9373922;
publickey_row[2732] = `CIPHERTEXT_WIDTH'd3637852;
publickey_row[2733] = `CIPHERTEXT_WIDTH'd452604;
publickey_row[2734] = `CIPHERTEXT_WIDTH'd7176227;
publickey_row[2735] = `CIPHERTEXT_WIDTH'd10135097;
publickey_row[2736] = `CIPHERTEXT_WIDTH'd11553856;
publickey_row[2737] = `CIPHERTEXT_WIDTH'd1690017;
publickey_row[2738] = `CIPHERTEXT_WIDTH'd5427869;
publickey_row[2739] = `CIPHERTEXT_WIDTH'd12902345;
publickey_row[2740] = `CIPHERTEXT_WIDTH'd4833197;
publickey_row[2741] = `CIPHERTEXT_WIDTH'd1498616;
publickey_row[2742] = `CIPHERTEXT_WIDTH'd7062682;
publickey_row[2743] = `CIPHERTEXT_WIDTH'd7039750;
publickey_row[2744] = `CIPHERTEXT_WIDTH'd1520317;
publickey_row[2745] = `CIPHERTEXT_WIDTH'd16270269;
publickey_row[2746] = `CIPHERTEXT_WIDTH'd12532896;
publickey_row[2747] = `CIPHERTEXT_WIDTH'd14813565;
publickey_row[2748] = `CIPHERTEXT_WIDTH'd12328929;
publickey_row[2749] = `CIPHERTEXT_WIDTH'd14206147;
publickey_row[2750] = `CIPHERTEXT_WIDTH'd14454996;
publickey_row[2751] = `CIPHERTEXT_WIDTH'd11646257;
publickey_row[2752] = `CIPHERTEXT_WIDTH'd4128710;
publickey_row[2753] = `CIPHERTEXT_WIDTH'd9367403;
publickey_row[2754] = `CIPHERTEXT_WIDTH'd6325377;
publickey_row[2755] = `CIPHERTEXT_WIDTH'd782086;
publickey_row[2756] = `CIPHERTEXT_WIDTH'd11214573;
publickey_row[2757] = `CIPHERTEXT_WIDTH'd10537157;
publickey_row[2758] = `CIPHERTEXT_WIDTH'd12728938;
publickey_row[2759] = `CIPHERTEXT_WIDTH'd16048923;
publickey_row[2760] = `CIPHERTEXT_WIDTH'd5603256;
publickey_row[2761] = `CIPHERTEXT_WIDTH'd4748300;
publickey_row[2762] = `CIPHERTEXT_WIDTH'd3584011;
publickey_row[2763] = `CIPHERTEXT_WIDTH'd7849430;
publickey_row[2764] = `CIPHERTEXT_WIDTH'd5542225;
publickey_row[2765] = `CIPHERTEXT_WIDTH'd7939244;
publickey_row[2766] = `CIPHERTEXT_WIDTH'd11022464;
publickey_row[2767] = `CIPHERTEXT_WIDTH'd164248;
publickey_row[2768] = `CIPHERTEXT_WIDTH'd14864686;
publickey_row[2769] = `CIPHERTEXT_WIDTH'd14494401;
publickey_row[2770] = `CIPHERTEXT_WIDTH'd450576;
publickey_row[2771] = `CIPHERTEXT_WIDTH'd11504323;
publickey_row[2772] = `CIPHERTEXT_WIDTH'd13553807;
publickey_row[2773] = `CIPHERTEXT_WIDTH'd896100;
publickey_row[2774] = `CIPHERTEXT_WIDTH'd3352508;
publickey_row[2775] = `CIPHERTEXT_WIDTH'd5998792;
publickey_row[2776] = `CIPHERTEXT_WIDTH'd8426681;
publickey_row[2777] = `CIPHERTEXT_WIDTH'd8149991;
publickey_row[2778] = `CIPHERTEXT_WIDTH'd3156559;
publickey_row[2779] = `CIPHERTEXT_WIDTH'd14318335;
publickey_row[2780] = `CIPHERTEXT_WIDTH'd8510859;
publickey_row[2781] = `CIPHERTEXT_WIDTH'd858235;
publickey_row[2782] = `CIPHERTEXT_WIDTH'd3795665;
publickey_row[2783] = `CIPHERTEXT_WIDTH'd12332068;
publickey_row[2784] = `CIPHERTEXT_WIDTH'd15939524;
publickey_row[2785] = `CIPHERTEXT_WIDTH'd6542325;
publickey_row[2786] = `CIPHERTEXT_WIDTH'd8271234;
publickey_row[2787] = `CIPHERTEXT_WIDTH'd9884897;
publickey_row[2788] = `CIPHERTEXT_WIDTH'd14840334;
publickey_row[2789] = `CIPHERTEXT_WIDTH'd641445;
publickey_row[2790] = `CIPHERTEXT_WIDTH'd15519730;
publickey_row[2791] = `CIPHERTEXT_WIDTH'd5432370;
publickey_row[2792] = `CIPHERTEXT_WIDTH'd6566110;
publickey_row[2793] = `CIPHERTEXT_WIDTH'd12396878;
publickey_row[2794] = `CIPHERTEXT_WIDTH'd15544316;
publickey_row[2795] = `CIPHERTEXT_WIDTH'd740293;
publickey_row[2796] = `CIPHERTEXT_WIDTH'd10746791;
publickey_row[2797] = `CIPHERTEXT_WIDTH'd6471411;
publickey_row[2798] = `CIPHERTEXT_WIDTH'd12809595;
publickey_row[2799] = `CIPHERTEXT_WIDTH'd8748090;
publickey_row[2800] = `CIPHERTEXT_WIDTH'd9290991;
publickey_row[2801] = `CIPHERTEXT_WIDTH'd3637460;
publickey_row[2802] = `CIPHERTEXT_WIDTH'd8842386;
publickey_row[2803] = `CIPHERTEXT_WIDTH'd9909702;
publickey_row[2804] = `CIPHERTEXT_WIDTH'd3371881;
publickey_row[2805] = `CIPHERTEXT_WIDTH'd3647327;
publickey_row[2806] = `CIPHERTEXT_WIDTH'd12432670;
publickey_row[2807] = `CIPHERTEXT_WIDTH'd1212828;
publickey_row[2808] = `CIPHERTEXT_WIDTH'd13915687;
publickey_row[2809] = `CIPHERTEXT_WIDTH'd14041090;
publickey_row[2810] = `CIPHERTEXT_WIDTH'd6039841;
publickey_row[2811] = `CIPHERTEXT_WIDTH'd5145219;
publickey_row[2812] = `CIPHERTEXT_WIDTH'd5884294;
publickey_row[2813] = `CIPHERTEXT_WIDTH'd8895483;
publickey_row[2814] = `CIPHERTEXT_WIDTH'd13171832;
publickey_row[2815] = `CIPHERTEXT_WIDTH'd3453998;
publickey_row[2816] = `CIPHERTEXT_WIDTH'd9555079;
publickey_row[2817] = `CIPHERTEXT_WIDTH'd1065130;
publickey_row[2818] = `CIPHERTEXT_WIDTH'd7317445;
publickey_row[2819] = `CIPHERTEXT_WIDTH'd8044483;
publickey_row[2820] = `CIPHERTEXT_WIDTH'd2835046;
publickey_row[2821] = `CIPHERTEXT_WIDTH'd6289454;
publickey_row[2822] = `CIPHERTEXT_WIDTH'd1910830;
publickey_row[2823] = `CIPHERTEXT_WIDTH'd15665296;
publickey_row[2824] = `CIPHERTEXT_WIDTH'd6680129;
publickey_row[2825] = `CIPHERTEXT_WIDTH'd16106011;
publickey_row[2826] = `CIPHERTEXT_WIDTH'd11228838;
publickey_row[2827] = `CIPHERTEXT_WIDTH'd564374;
publickey_row[2828] = `CIPHERTEXT_WIDTH'd13400702;
publickey_row[2829] = `CIPHERTEXT_WIDTH'd10959779;
publickey_row[2830] = `CIPHERTEXT_WIDTH'd64667;
publickey_row[2831] = `CIPHERTEXT_WIDTH'd4432466;
publickey_row[2832] = `CIPHERTEXT_WIDTH'd6960798;
publickey_row[2833] = `CIPHERTEXT_WIDTH'd4273538;
publickey_row[2834] = `CIPHERTEXT_WIDTH'd8424207;
publickey_row[2835] = `CIPHERTEXT_WIDTH'd3815164;
publickey_row[2836] = `CIPHERTEXT_WIDTH'd822885;
publickey_row[2837] = `CIPHERTEXT_WIDTH'd16396005;
publickey_row[2838] = `CIPHERTEXT_WIDTH'd10408812;
publickey_row[2839] = `CIPHERTEXT_WIDTH'd8445416;
publickey_row[2840] = `CIPHERTEXT_WIDTH'd70814;
publickey_row[2841] = `CIPHERTEXT_WIDTH'd13126753;
publickey_row[2842] = `CIPHERTEXT_WIDTH'd4667708;
publickey_row[2843] = `CIPHERTEXT_WIDTH'd9429062;
publickey_row[2844] = `CIPHERTEXT_WIDTH'd1888731;
publickey_row[2845] = `CIPHERTEXT_WIDTH'd13836408;
publickey_row[2846] = `CIPHERTEXT_WIDTH'd1417195;
publickey_row[2847] = `CIPHERTEXT_WIDTH'd10496393;
publickey_row[2848] = `CIPHERTEXT_WIDTH'd6010190;
publickey_row[2849] = `CIPHERTEXT_WIDTH'd7985682;
publickey_row[2850] = `CIPHERTEXT_WIDTH'd13898416;
publickey_row[2851] = `CIPHERTEXT_WIDTH'd11512126;
publickey_row[2852] = `CIPHERTEXT_WIDTH'd5650861;
publickey_row[2853] = `CIPHERTEXT_WIDTH'd12408329;
publickey_row[2854] = `CIPHERTEXT_WIDTH'd16671776;
publickey_row[2855] = `CIPHERTEXT_WIDTH'd3122307;
publickey_row[2856] = `CIPHERTEXT_WIDTH'd9150368;
publickey_row[2857] = `CIPHERTEXT_WIDTH'd8762950;
publickey_row[2858] = `CIPHERTEXT_WIDTH'd1843681;
publickey_row[2859] = `CIPHERTEXT_WIDTH'd14310685;
publickey_row[2860] = `CIPHERTEXT_WIDTH'd12744779;
publickey_row[2861] = `CIPHERTEXT_WIDTH'd10544379;
publickey_row[2862] = `CIPHERTEXT_WIDTH'd2735459;
publickey_row[2863] = `CIPHERTEXT_WIDTH'd2893952;
publickey_row[2864] = `CIPHERTEXT_WIDTH'd14709410;
publickey_row[2865] = `CIPHERTEXT_WIDTH'd948314;
publickey_row[2866] = `CIPHERTEXT_WIDTH'd2441400;
publickey_row[2867] = `CIPHERTEXT_WIDTH'd14995948;
publickey_row[2868] = `CIPHERTEXT_WIDTH'd3478011;
publickey_row[2869] = `CIPHERTEXT_WIDTH'd606273;
publickey_row[2870] = `CIPHERTEXT_WIDTH'd15414273;
publickey_row[2871] = `CIPHERTEXT_WIDTH'd14438173;
publickey_row[2872] = `CIPHERTEXT_WIDTH'd13178109;
publickey_row[2873] = `CIPHERTEXT_WIDTH'd7296498;
publickey_row[2874] = `CIPHERTEXT_WIDTH'd3827696;
publickey_row[2875] = `CIPHERTEXT_WIDTH'd11459285;
publickey_row[2876] = `CIPHERTEXT_WIDTH'd11110559;
publickey_row[2877] = `CIPHERTEXT_WIDTH'd15819688;
publickey_row[2878] = `CIPHERTEXT_WIDTH'd6585375;
publickey_row[2879] = `CIPHERTEXT_WIDTH'd5635959;
publickey_row[2880] = `CIPHERTEXT_WIDTH'd15942007;
publickey_row[2881] = `CIPHERTEXT_WIDTH'd8953155;
publickey_row[2882] = `CIPHERTEXT_WIDTH'd1247044;
publickey_row[2883] = `CIPHERTEXT_WIDTH'd5658020;
publickey_row[2884] = `CIPHERTEXT_WIDTH'd14894252;
publickey_row[2885] = `CIPHERTEXT_WIDTH'd444095;
publickey_row[2886] = `CIPHERTEXT_WIDTH'd975395;
publickey_row[2887] = `CIPHERTEXT_WIDTH'd16275386;
publickey_row[2888] = `CIPHERTEXT_WIDTH'd550882;
publickey_row[2889] = `CIPHERTEXT_WIDTH'd438786;
publickey_row[2890] = `CIPHERTEXT_WIDTH'd15360361;
publickey_row[2891] = `CIPHERTEXT_WIDTH'd14626355;
publickey_row[2892] = `CIPHERTEXT_WIDTH'd14979098;
publickey_row[2893] = `CIPHERTEXT_WIDTH'd286057;
publickey_row[2894] = `CIPHERTEXT_WIDTH'd4926058;
publickey_row[2895] = `CIPHERTEXT_WIDTH'd11364290;
publickey_row[2896] = `CIPHERTEXT_WIDTH'd16676795;
publickey_row[2897] = `CIPHERTEXT_WIDTH'd15514446;
publickey_row[2898] = `CIPHERTEXT_WIDTH'd4116371;
publickey_row[2899] = `CIPHERTEXT_WIDTH'd13436135;
publickey_row[2900] = `CIPHERTEXT_WIDTH'd13222368;
publickey_row[2901] = `CIPHERTEXT_WIDTH'd11215035;
publickey_row[2902] = `CIPHERTEXT_WIDTH'd1104008;
publickey_row[2903] = `CIPHERTEXT_WIDTH'd561452;
publickey_row[2904] = `CIPHERTEXT_WIDTH'd1648299;
publickey_row[2905] = `CIPHERTEXT_WIDTH'd6025964;
publickey_row[2906] = `CIPHERTEXT_WIDTH'd5585995;
publickey_row[2907] = `CIPHERTEXT_WIDTH'd10354414;
publickey_row[2908] = `CIPHERTEXT_WIDTH'd5143704;
publickey_row[2909] = `CIPHERTEXT_WIDTH'd1282922;
publickey_row[2910] = `CIPHERTEXT_WIDTH'd12828608;
publickey_row[2911] = `CIPHERTEXT_WIDTH'd12773741;
publickey_row[2912] = `CIPHERTEXT_WIDTH'd15848573;
publickey_row[2913] = `CIPHERTEXT_WIDTH'd188464;
publickey_row[2914] = `CIPHERTEXT_WIDTH'd5265121;
publickey_row[2915] = `CIPHERTEXT_WIDTH'd7771608;
publickey_row[2916] = `CIPHERTEXT_WIDTH'd5818158;
publickey_row[2917] = `CIPHERTEXT_WIDTH'd12361700;
publickey_row[2918] = `CIPHERTEXT_WIDTH'd11812997;
publickey_row[2919] = `CIPHERTEXT_WIDTH'd9617198;
publickey_row[2920] = `CIPHERTEXT_WIDTH'd15031168;
publickey_row[2921] = `CIPHERTEXT_WIDTH'd7731302;
publickey_row[2922] = `CIPHERTEXT_WIDTH'd10288842;
publickey_row[2923] = `CIPHERTEXT_WIDTH'd12208761;
publickey_row[2924] = `CIPHERTEXT_WIDTH'd5484228;
publickey_row[2925] = `CIPHERTEXT_WIDTH'd3178678;
publickey_row[2926] = `CIPHERTEXT_WIDTH'd7339743;
publickey_row[2927] = `CIPHERTEXT_WIDTH'd9546339;
publickey_row[2928] = `CIPHERTEXT_WIDTH'd16700481;
publickey_row[2929] = `CIPHERTEXT_WIDTH'd3064297;
publickey_row[2930] = `CIPHERTEXT_WIDTH'd9699091;
publickey_row[2931] = `CIPHERTEXT_WIDTH'd15255386;
publickey_row[2932] = `CIPHERTEXT_WIDTH'd6467987;
publickey_row[2933] = `CIPHERTEXT_WIDTH'd15389240;
publickey_row[2934] = `CIPHERTEXT_WIDTH'd936525;
publickey_row[2935] = `CIPHERTEXT_WIDTH'd4679047;
publickey_row[2936] = `CIPHERTEXT_WIDTH'd9171304;
publickey_row[2937] = `CIPHERTEXT_WIDTH'd10026453;
publickey_row[2938] = `CIPHERTEXT_WIDTH'd12318030;
publickey_row[2939] = `CIPHERTEXT_WIDTH'd9157160;
publickey_row[2940] = `CIPHERTEXT_WIDTH'd11634123;
publickey_row[2941] = `CIPHERTEXT_WIDTH'd3304419;
publickey_row[2942] = `CIPHERTEXT_WIDTH'd1476486;
publickey_row[2943] = `CIPHERTEXT_WIDTH'd13487644;
publickey_row[2944] = `CIPHERTEXT_WIDTH'd13735554;
publickey_row[2945] = `CIPHERTEXT_WIDTH'd10613495;
publickey_row[2946] = `CIPHERTEXT_WIDTH'd14808410;
publickey_row[2947] = `CIPHERTEXT_WIDTH'd5443018;
publickey_row[2948] = `CIPHERTEXT_WIDTH'd1005970;
publickey_row[2949] = `CIPHERTEXT_WIDTH'd5635882;
publickey_row[2950] = `CIPHERTEXT_WIDTH'd15759197;
publickey_row[2951] = `CIPHERTEXT_WIDTH'd15314889;
publickey_row[2952] = `CIPHERTEXT_WIDTH'd2186741;
publickey_row[2953] = `CIPHERTEXT_WIDTH'd14686776;
publickey_row[2954] = `CIPHERTEXT_WIDTH'd927576;
publickey_row[2955] = `CIPHERTEXT_WIDTH'd6309355;
publickey_row[2956] = `CIPHERTEXT_WIDTH'd8357965;
publickey_row[2957] = `CIPHERTEXT_WIDTH'd13852446;
publickey_row[2958] = `CIPHERTEXT_WIDTH'd3096689;
publickey_row[2959] = `CIPHERTEXT_WIDTH'd94295;
publickey_row[2960] = `CIPHERTEXT_WIDTH'd13018084;
publickey_row[2961] = `CIPHERTEXT_WIDTH'd5599608;
publickey_row[2962] = `CIPHERTEXT_WIDTH'd16675021;
publickey_row[2963] = `CIPHERTEXT_WIDTH'd13952588;
publickey_row[2964] = `CIPHERTEXT_WIDTH'd16729306;
publickey_row[2965] = `CIPHERTEXT_WIDTH'd15611674;
publickey_row[2966] = `CIPHERTEXT_WIDTH'd6834914;
publickey_row[2967] = `CIPHERTEXT_WIDTH'd1665670;
publickey_row[2968] = `CIPHERTEXT_WIDTH'd10854395;
publickey_row[2969] = `CIPHERTEXT_WIDTH'd10538973;
publickey_row[2970] = `CIPHERTEXT_WIDTH'd9134332;
publickey_row[2971] = `CIPHERTEXT_WIDTH'd12093123;
publickey_row[2972] = `CIPHERTEXT_WIDTH'd14179885;
publickey_row[2973] = `CIPHERTEXT_WIDTH'd15829972;
publickey_row[2974] = `CIPHERTEXT_WIDTH'd974515;
publickey_row[2975] = `CIPHERTEXT_WIDTH'd927164;
publickey_row[2976] = `CIPHERTEXT_WIDTH'd7064396;
publickey_row[2977] = `CIPHERTEXT_WIDTH'd6110394;
publickey_row[2978] = `CIPHERTEXT_WIDTH'd11520452;
publickey_row[2979] = `CIPHERTEXT_WIDTH'd13468710;
publickey_row[2980] = `CIPHERTEXT_WIDTH'd13763640;
publickey_row[2981] = `CIPHERTEXT_WIDTH'd5401627;
publickey_row[2982] = `CIPHERTEXT_WIDTH'd15929002;
publickey_row[2983] = `CIPHERTEXT_WIDTH'd11641845;
publickey_row[2984] = `CIPHERTEXT_WIDTH'd4139639;
publickey_row[2985] = `CIPHERTEXT_WIDTH'd1960517;
publickey_row[2986] = `CIPHERTEXT_WIDTH'd11480537;
publickey_row[2987] = `CIPHERTEXT_WIDTH'd1713504;
publickey_row[2988] = `CIPHERTEXT_WIDTH'd12063243;
publickey_row[2989] = `CIPHERTEXT_WIDTH'd11403193;
publickey_row[2990] = `CIPHERTEXT_WIDTH'd7191388;
publickey_row[2991] = `CIPHERTEXT_WIDTH'd13011810;
publickey_row[2992] = `CIPHERTEXT_WIDTH'd16691113;
publickey_row[2993] = `CIPHERTEXT_WIDTH'd6943280;
publickey_row[2994] = `CIPHERTEXT_WIDTH'd4991193;
publickey_row[2995] = `CIPHERTEXT_WIDTH'd3151767;
publickey_row[2996] = `CIPHERTEXT_WIDTH'd519134;
publickey_row[2997] = `CIPHERTEXT_WIDTH'd14723043;
publickey_row[2998] = `CIPHERTEXT_WIDTH'd9904466;
publickey_row[2999] = `CIPHERTEXT_WIDTH'd12736202;
publickey_row[3000] = `CIPHERTEXT_WIDTH'd11361043;
publickey_row[3001] = `CIPHERTEXT_WIDTH'd5394851;
publickey_row[3002] = `CIPHERTEXT_WIDTH'd5268878;
publickey_row[3003] = `CIPHERTEXT_WIDTH'd15971243;
publickey_row[3004] = `CIPHERTEXT_WIDTH'd16103843;
publickey_row[3005] = `CIPHERTEXT_WIDTH'd283357;
publickey_row[3006] = `CIPHERTEXT_WIDTH'd857246;
publickey_row[3007] = `CIPHERTEXT_WIDTH'd1361053;
publickey_row[3008] = `CIPHERTEXT_WIDTH'd4194523;
publickey_row[3009] = `CIPHERTEXT_WIDTH'd4288476;
publickey_row[3010] = `CIPHERTEXT_WIDTH'd5642759;
publickey_row[3011] = `CIPHERTEXT_WIDTH'd4470316;
publickey_row[3012] = `CIPHERTEXT_WIDTH'd7868982;
publickey_row[3013] = `CIPHERTEXT_WIDTH'd15449634;
publickey_row[3014] = `CIPHERTEXT_WIDTH'd624886;
publickey_row[3015] = `CIPHERTEXT_WIDTH'd1689761;
publickey_row[3016] = `CIPHERTEXT_WIDTH'd2773295;
publickey_row[3017] = `CIPHERTEXT_WIDTH'd4769054;
publickey_row[3018] = `CIPHERTEXT_WIDTH'd10366717;
publickey_row[3019] = `CIPHERTEXT_WIDTH'd2555159;
publickey_row[3020] = `CIPHERTEXT_WIDTH'd5544844;
publickey_row[3021] = `CIPHERTEXT_WIDTH'd4309132;
publickey_row[3022] = `CIPHERTEXT_WIDTH'd11145018;
publickey_row[3023] = `CIPHERTEXT_WIDTH'd12594884;
publickey_row[3024] = `CIPHERTEXT_WIDTH'd15460947;
publickey_row[3025] = `CIPHERTEXT_WIDTH'd5518757;
publickey_row[3026] = `CIPHERTEXT_WIDTH'd3328240;
publickey_row[3027] = `CIPHERTEXT_WIDTH'd1931171;
publickey_row[3028] = `CIPHERTEXT_WIDTH'd5380435;
publickey_row[3029] = `CIPHERTEXT_WIDTH'd11856344;
publickey_row[3030] = `CIPHERTEXT_WIDTH'd12741815;
publickey_row[3031] = `CIPHERTEXT_WIDTH'd8746498;
publickey_row[3032] = `CIPHERTEXT_WIDTH'd15196168;
publickey_row[3033] = `CIPHERTEXT_WIDTH'd11373754;
publickey_row[3034] = `CIPHERTEXT_WIDTH'd13927252;
publickey_row[3035] = `CIPHERTEXT_WIDTH'd6106036;
publickey_row[3036] = `CIPHERTEXT_WIDTH'd957223;
publickey_row[3037] = `CIPHERTEXT_WIDTH'd8193323;
publickey_row[3038] = `CIPHERTEXT_WIDTH'd12410425;
publickey_row[3039] = `CIPHERTEXT_WIDTH'd9880681;
publickey_row[3040] = `CIPHERTEXT_WIDTH'd1904556;
publickey_row[3041] = `CIPHERTEXT_WIDTH'd2859813;
publickey_row[3042] = `CIPHERTEXT_WIDTH'd16689704;
publickey_row[3043] = `CIPHERTEXT_WIDTH'd16584246;
publickey_row[3044] = `CIPHERTEXT_WIDTH'd2409432;
publickey_row[3045] = `CIPHERTEXT_WIDTH'd14696097;
publickey_row[3046] = `CIPHERTEXT_WIDTH'd13528413;
publickey_row[3047] = `CIPHERTEXT_WIDTH'd10116223;
publickey_row[3048] = `CIPHERTEXT_WIDTH'd9078072;
publickey_row[3049] = `CIPHERTEXT_WIDTH'd15133212;
publickey_row[3050] = `CIPHERTEXT_WIDTH'd10887836;
publickey_row[3051] = `CIPHERTEXT_WIDTH'd9693889;
publickey_row[3052] = `CIPHERTEXT_WIDTH'd14056863;
publickey_row[3053] = `CIPHERTEXT_WIDTH'd3004870;
publickey_row[3054] = `CIPHERTEXT_WIDTH'd12234517;
publickey_row[3055] = `CIPHERTEXT_WIDTH'd14467711;
publickey_row[3056] = `CIPHERTEXT_WIDTH'd14740014;
publickey_row[3057] = `CIPHERTEXT_WIDTH'd6977049;
publickey_row[3058] = `CIPHERTEXT_WIDTH'd10518550;
publickey_row[3059] = `CIPHERTEXT_WIDTH'd14237856;
publickey_row[3060] = `CIPHERTEXT_WIDTH'd8249006;
publickey_row[3061] = `CIPHERTEXT_WIDTH'd12882292;
publickey_row[3062] = `CIPHERTEXT_WIDTH'd88131;
publickey_row[3063] = `CIPHERTEXT_WIDTH'd15657800;
publickey_row[3064] = `CIPHERTEXT_WIDTH'd13892956;
publickey_row[3065] = `CIPHERTEXT_WIDTH'd4769473;
publickey_row[3066] = `CIPHERTEXT_WIDTH'd15518400;
publickey_row[3067] = `CIPHERTEXT_WIDTH'd5469803;
publickey_row[3068] = `CIPHERTEXT_WIDTH'd6464128;
publickey_row[3069] = `CIPHERTEXT_WIDTH'd4072986;
publickey_row[3070] = `CIPHERTEXT_WIDTH'd15277938;
publickey_row[3071] = `CIPHERTEXT_WIDTH'd4657175;
publickey_row[3072] = `CIPHERTEXT_WIDTH'd6265877;
publickey_row[3073] = `CIPHERTEXT_WIDTH'd6734038;
publickey_row[3074] = `CIPHERTEXT_WIDTH'd3269827;
publickey_row[3075] = `CIPHERTEXT_WIDTH'd8507202;
publickey_row[3076] = `CIPHERTEXT_WIDTH'd10340567;
publickey_row[3077] = `CIPHERTEXT_WIDTH'd6173739;
publickey_row[3078] = `CIPHERTEXT_WIDTH'd13564756;
publickey_row[3079] = `CIPHERTEXT_WIDTH'd5811571;
publickey_row[3080] = `CIPHERTEXT_WIDTH'd2593772;
publickey_row[3081] = `CIPHERTEXT_WIDTH'd10171706;
publickey_row[3082] = `CIPHERTEXT_WIDTH'd12211372;
publickey_row[3083] = `CIPHERTEXT_WIDTH'd7274579;
publickey_row[3084] = `CIPHERTEXT_WIDTH'd1716204;
publickey_row[3085] = `CIPHERTEXT_WIDTH'd9868623;
publickey_row[3086] = `CIPHERTEXT_WIDTH'd5915983;
publickey_row[3087] = `CIPHERTEXT_WIDTH'd11335179;
publickey_row[3088] = `CIPHERTEXT_WIDTH'd12383054;
publickey_row[3089] = `CIPHERTEXT_WIDTH'd12167176;
publickey_row[3090] = `CIPHERTEXT_WIDTH'd364357;
publickey_row[3091] = `CIPHERTEXT_WIDTH'd2556976;
publickey_row[3092] = `CIPHERTEXT_WIDTH'd10658848;
publickey_row[3093] = `CIPHERTEXT_WIDTH'd23491;
publickey_row[3094] = `CIPHERTEXT_WIDTH'd5689693;
publickey_row[3095] = `CIPHERTEXT_WIDTH'd7233871;
publickey_row[3096] = `CIPHERTEXT_WIDTH'd16349054;
publickey_row[3097] = `CIPHERTEXT_WIDTH'd476595;
publickey_row[3098] = `CIPHERTEXT_WIDTH'd9150242;
publickey_row[3099] = `CIPHERTEXT_WIDTH'd4120983;
publickey_row[3100] = `CIPHERTEXT_WIDTH'd2828729;
publickey_row[3101] = `CIPHERTEXT_WIDTH'd8624745;
publickey_row[3102] = `CIPHERTEXT_WIDTH'd1336504;
publickey_row[3103] = `CIPHERTEXT_WIDTH'd11771597;
publickey_row[3104] = `CIPHERTEXT_WIDTH'd304495;
publickey_row[3105] = `CIPHERTEXT_WIDTH'd15615679;
publickey_row[3106] = `CIPHERTEXT_WIDTH'd6330141;
publickey_row[3107] = `CIPHERTEXT_WIDTH'd3272178;
publickey_row[3108] = `CIPHERTEXT_WIDTH'd9338023;
publickey_row[3109] = `CIPHERTEXT_WIDTH'd10871087;
publickey_row[3110] = `CIPHERTEXT_WIDTH'd11458312;
publickey_row[3111] = `CIPHERTEXT_WIDTH'd16458294;
publickey_row[3112] = `CIPHERTEXT_WIDTH'd14013179;
publickey_row[3113] = `CIPHERTEXT_WIDTH'd6245859;
publickey_row[3114] = `CIPHERTEXT_WIDTH'd2600616;
publickey_row[3115] = `CIPHERTEXT_WIDTH'd2020947;
publickey_row[3116] = `CIPHERTEXT_WIDTH'd7124118;
publickey_row[3117] = `CIPHERTEXT_WIDTH'd14954852;
publickey_row[3118] = `CIPHERTEXT_WIDTH'd1691456;
publickey_row[3119] = `CIPHERTEXT_WIDTH'd15224610;
publickey_row[3120] = `CIPHERTEXT_WIDTH'd15454409;
publickey_row[3121] = `CIPHERTEXT_WIDTH'd2265909;
publickey_row[3122] = `CIPHERTEXT_WIDTH'd876630;
publickey_row[3123] = `CIPHERTEXT_WIDTH'd2089781;
publickey_row[3124] = `CIPHERTEXT_WIDTH'd4631730;
publickey_row[3125] = `CIPHERTEXT_WIDTH'd6410176;
publickey_row[3126] = `CIPHERTEXT_WIDTH'd9726723;
publickey_row[3127] = `CIPHERTEXT_WIDTH'd12507671;
publickey_row[3128] = `CIPHERTEXT_WIDTH'd5070557;
publickey_row[3129] = `CIPHERTEXT_WIDTH'd13861829;
publickey_row[3130] = `CIPHERTEXT_WIDTH'd12989768;
publickey_row[3131] = `CIPHERTEXT_WIDTH'd11369915;
publickey_row[3132] = `CIPHERTEXT_WIDTH'd1559633;
publickey_row[3133] = `CIPHERTEXT_WIDTH'd8373672;
publickey_row[3134] = `CIPHERTEXT_WIDTH'd15487771;
publickey_row[3135] = `CIPHERTEXT_WIDTH'd1626344;
publickey_row[3136] = `CIPHERTEXT_WIDTH'd107852;
publickey_row[3137] = `CIPHERTEXT_WIDTH'd6009675;
publickey_row[3138] = `CIPHERTEXT_WIDTH'd6927872;
publickey_row[3139] = `CIPHERTEXT_WIDTH'd7969010;
publickey_row[3140] = `CIPHERTEXT_WIDTH'd3347643;
publickey_row[3141] = `CIPHERTEXT_WIDTH'd1424973;
publickey_row[3142] = `CIPHERTEXT_WIDTH'd2296608;
publickey_row[3143] = `CIPHERTEXT_WIDTH'd9022412;
publickey_row[3144] = `CIPHERTEXT_WIDTH'd9912117;
publickey_row[3145] = `CIPHERTEXT_WIDTH'd10166;
publickey_row[3146] = `CIPHERTEXT_WIDTH'd5392201;
publickey_row[3147] = `CIPHERTEXT_WIDTH'd4027225;
publickey_row[3148] = `CIPHERTEXT_WIDTH'd9885040;
publickey_row[3149] = `CIPHERTEXT_WIDTH'd16248402;
publickey_row[3150] = `CIPHERTEXT_WIDTH'd1664838;
publickey_row[3151] = `CIPHERTEXT_WIDTH'd5922913;
publickey_row[3152] = `CIPHERTEXT_WIDTH'd893188;
publickey_row[3153] = `CIPHERTEXT_WIDTH'd7967988;
publickey_row[3154] = `CIPHERTEXT_WIDTH'd6321301;
publickey_row[3155] = `CIPHERTEXT_WIDTH'd10383870;
publickey_row[3156] = `CIPHERTEXT_WIDTH'd10160830;
publickey_row[3157] = `CIPHERTEXT_WIDTH'd15939359;
publickey_row[3158] = `CIPHERTEXT_WIDTH'd4515320;
publickey_row[3159] = `CIPHERTEXT_WIDTH'd2866031;
publickey_row[3160] = `CIPHERTEXT_WIDTH'd15506510;
publickey_row[3161] = `CIPHERTEXT_WIDTH'd16759853;
publickey_row[3162] = `CIPHERTEXT_WIDTH'd15822108;
publickey_row[3163] = `CIPHERTEXT_WIDTH'd5804062;
publickey_row[3164] = `CIPHERTEXT_WIDTH'd12685828;
publickey_row[3165] = `CIPHERTEXT_WIDTH'd3982764;
publickey_row[3166] = `CIPHERTEXT_WIDTH'd8098258;
publickey_row[3167] = `CIPHERTEXT_WIDTH'd6425828;
publickey_row[3168] = `CIPHERTEXT_WIDTH'd3642638;
publickey_row[3169] = `CIPHERTEXT_WIDTH'd5660643;
publickey_row[3170] = `CIPHERTEXT_WIDTH'd15632528;
publickey_row[3171] = `CIPHERTEXT_WIDTH'd6795347;
publickey_row[3172] = `CIPHERTEXT_WIDTH'd10824126;
publickey_row[3173] = `CIPHERTEXT_WIDTH'd5607119;
publickey_row[3174] = `CIPHERTEXT_WIDTH'd13870119;
publickey_row[3175] = `CIPHERTEXT_WIDTH'd14305787;
publickey_row[3176] = `CIPHERTEXT_WIDTH'd2852692;
publickey_row[3177] = `CIPHERTEXT_WIDTH'd3930035;
publickey_row[3178] = `CIPHERTEXT_WIDTH'd732449;
publickey_row[3179] = `CIPHERTEXT_WIDTH'd2437261;
publickey_row[3180] = `CIPHERTEXT_WIDTH'd14908197;
publickey_row[3181] = `CIPHERTEXT_WIDTH'd14616624;
publickey_row[3182] = `CIPHERTEXT_WIDTH'd3343184;
publickey_row[3183] = `CIPHERTEXT_WIDTH'd8338007;
publickey_row[3184] = `CIPHERTEXT_WIDTH'd5993814;
publickey_row[3185] = `CIPHERTEXT_WIDTH'd5587517;
publickey_row[3186] = `CIPHERTEXT_WIDTH'd14393527;
publickey_row[3187] = `CIPHERTEXT_WIDTH'd1252267;
publickey_row[3188] = `CIPHERTEXT_WIDTH'd1460065;
publickey_row[3189] = `CIPHERTEXT_WIDTH'd2447878;
publickey_row[3190] = `CIPHERTEXT_WIDTH'd14204486;
publickey_row[3191] = `CIPHERTEXT_WIDTH'd659712;
publickey_row[3192] = `CIPHERTEXT_WIDTH'd6275186;
publickey_row[3193] = `CIPHERTEXT_WIDTH'd557163;
publickey_row[3194] = `CIPHERTEXT_WIDTH'd69188;
publickey_row[3195] = `CIPHERTEXT_WIDTH'd5401949;
publickey_row[3196] = `CIPHERTEXT_WIDTH'd5176790;
publickey_row[3197] = `CIPHERTEXT_WIDTH'd5696665;
publickey_row[3198] = `CIPHERTEXT_WIDTH'd14423294;
publickey_row[3199] = `CIPHERTEXT_WIDTH'd9349310;
publickey_row[3200] = `CIPHERTEXT_WIDTH'd16519836;
publickey_row[3201] = `CIPHERTEXT_WIDTH'd16352591;
publickey_row[3202] = `CIPHERTEXT_WIDTH'd12000472;
publickey_row[3203] = `CIPHERTEXT_WIDTH'd5471552;
publickey_row[3204] = `CIPHERTEXT_WIDTH'd5157978;
publickey_row[3205] = `CIPHERTEXT_WIDTH'd2482413;
publickey_row[3206] = `CIPHERTEXT_WIDTH'd2612390;
publickey_row[3207] = `CIPHERTEXT_WIDTH'd476254;
publickey_row[3208] = `CIPHERTEXT_WIDTH'd6960533;
publickey_row[3209] = `CIPHERTEXT_WIDTH'd935714;
publickey_row[3210] = `CIPHERTEXT_WIDTH'd14425541;
publickey_row[3211] = `CIPHERTEXT_WIDTH'd4584168;
publickey_row[3212] = `CIPHERTEXT_WIDTH'd12023511;
publickey_row[3213] = `CIPHERTEXT_WIDTH'd472511;
publickey_row[3214] = `CIPHERTEXT_WIDTH'd6961937;
publickey_row[3215] = `CIPHERTEXT_WIDTH'd2492610;
publickey_row[3216] = `CIPHERTEXT_WIDTH'd3037698;
publickey_row[3217] = `CIPHERTEXT_WIDTH'd751707;
publickey_row[3218] = `CIPHERTEXT_WIDTH'd2180324;
publickey_row[3219] = `CIPHERTEXT_WIDTH'd1542553;
publickey_row[3220] = `CIPHERTEXT_WIDTH'd15850879;
publickey_row[3221] = `CIPHERTEXT_WIDTH'd2766093;
publickey_row[3222] = `CIPHERTEXT_WIDTH'd442369;
publickey_row[3223] = `CIPHERTEXT_WIDTH'd8932818;
publickey_row[3224] = `CIPHERTEXT_WIDTH'd11375583;
publickey_row[3225] = `CIPHERTEXT_WIDTH'd12066255;
publickey_row[3226] = `CIPHERTEXT_WIDTH'd8680849;
publickey_row[3227] = `CIPHERTEXT_WIDTH'd15707089;
publickey_row[3228] = `CIPHERTEXT_WIDTH'd12250889;
publickey_row[3229] = `CIPHERTEXT_WIDTH'd4553958;
publickey_row[3230] = `CIPHERTEXT_WIDTH'd6710578;
publickey_row[3231] = `CIPHERTEXT_WIDTH'd16238597;
publickey_row[3232] = `CIPHERTEXT_WIDTH'd15326360;
publickey_row[3233] = `CIPHERTEXT_WIDTH'd3951331;
publickey_row[3234] = `CIPHERTEXT_WIDTH'd9704290;
publickey_row[3235] = `CIPHERTEXT_WIDTH'd820269;
publickey_row[3236] = `CIPHERTEXT_WIDTH'd7779216;
publickey_row[3237] = `CIPHERTEXT_WIDTH'd12204157;
publickey_row[3238] = `CIPHERTEXT_WIDTH'd12723851;
publickey_row[3239] = `CIPHERTEXT_WIDTH'd14872095;
publickey_row[3240] = `CIPHERTEXT_WIDTH'd11316833;
publickey_row[3241] = `CIPHERTEXT_WIDTH'd80997;
publickey_row[3242] = `CIPHERTEXT_WIDTH'd4328054;
publickey_row[3243] = `CIPHERTEXT_WIDTH'd1658071;
publickey_row[3244] = `CIPHERTEXT_WIDTH'd10630835;
publickey_row[3245] = `CIPHERTEXT_WIDTH'd15186350;
publickey_row[3246] = `CIPHERTEXT_WIDTH'd1177869;
publickey_row[3247] = `CIPHERTEXT_WIDTH'd3611456;
publickey_row[3248] = `CIPHERTEXT_WIDTH'd9021328;
publickey_row[3249] = `CIPHERTEXT_WIDTH'd4327878;
publickey_row[3250] = `CIPHERTEXT_WIDTH'd12377908;
publickey_row[3251] = `CIPHERTEXT_WIDTH'd16256600;
publickey_row[3252] = `CIPHERTEXT_WIDTH'd3644496;
publickey_row[3253] = `CIPHERTEXT_WIDTH'd5546064;
publickey_row[3254] = `CIPHERTEXT_WIDTH'd2108194;
publickey_row[3255] = `CIPHERTEXT_WIDTH'd14121794;
publickey_row[3256] = `CIPHERTEXT_WIDTH'd10425232;
publickey_row[3257] = `CIPHERTEXT_WIDTH'd4388552;
publickey_row[3258] = `CIPHERTEXT_WIDTH'd14819709;
publickey_row[3259] = `CIPHERTEXT_WIDTH'd5192501;
publickey_row[3260] = `CIPHERTEXT_WIDTH'd12167693;
publickey_row[3261] = `CIPHERTEXT_WIDTH'd14081330;
publickey_row[3262] = `CIPHERTEXT_WIDTH'd12749581;
publickey_row[3263] = `CIPHERTEXT_WIDTH'd4624618;
publickey_row[3264] = `CIPHERTEXT_WIDTH'd7191602;
publickey_row[3265] = `CIPHERTEXT_WIDTH'd7762493;
publickey_row[3266] = `CIPHERTEXT_WIDTH'd5005013;
publickey_row[3267] = `CIPHERTEXT_WIDTH'd60920;
publickey_row[3268] = `CIPHERTEXT_WIDTH'd8420090;
publickey_row[3269] = `CIPHERTEXT_WIDTH'd11709540;
publickey_row[3270] = `CIPHERTEXT_WIDTH'd4739972;
publickey_row[3271] = `CIPHERTEXT_WIDTH'd7346165;
publickey_row[3272] = `CIPHERTEXT_WIDTH'd5306875;
publickey_row[3273] = `CIPHERTEXT_WIDTH'd13990564;
publickey_row[3274] = `CIPHERTEXT_WIDTH'd7827575;
publickey_row[3275] = `CIPHERTEXT_WIDTH'd9431963;
publickey_row[3276] = `CIPHERTEXT_WIDTH'd5552083;
publickey_row[3277] = `CIPHERTEXT_WIDTH'd3264438;
publickey_row[3278] = `CIPHERTEXT_WIDTH'd4854109;
publickey_row[3279] = `CIPHERTEXT_WIDTH'd4527220;
publickey_row[3280] = `CIPHERTEXT_WIDTH'd12090020;
publickey_row[3281] = `CIPHERTEXT_WIDTH'd14476448;
publickey_row[3282] = `CIPHERTEXT_WIDTH'd7305004;
publickey_row[3283] = `CIPHERTEXT_WIDTH'd4718935;
publickey_row[3284] = `CIPHERTEXT_WIDTH'd6681938;
publickey_row[3285] = `CIPHERTEXT_WIDTH'd9681175;
publickey_row[3286] = `CIPHERTEXT_WIDTH'd6842426;
publickey_row[3287] = `CIPHERTEXT_WIDTH'd13613743;
publickey_row[3288] = `CIPHERTEXT_WIDTH'd11991443;
publickey_row[3289] = `CIPHERTEXT_WIDTH'd11884842;
publickey_row[3290] = `CIPHERTEXT_WIDTH'd429282;
publickey_row[3291] = `CIPHERTEXT_WIDTH'd3585639;
publickey_row[3292] = `CIPHERTEXT_WIDTH'd313997;
publickey_row[3293] = `CIPHERTEXT_WIDTH'd8381808;
publickey_row[3294] = `CIPHERTEXT_WIDTH'd6406317;
publickey_row[3295] = `CIPHERTEXT_WIDTH'd9951537;
publickey_row[3296] = `CIPHERTEXT_WIDTH'd6819100;
publickey_row[3297] = `CIPHERTEXT_WIDTH'd15280050;
publickey_row[3298] = `CIPHERTEXT_WIDTH'd12732463;
publickey_row[3299] = `CIPHERTEXT_WIDTH'd7837421;
publickey_row[3300] = `CIPHERTEXT_WIDTH'd14719333;
publickey_row[3301] = `CIPHERTEXT_WIDTH'd6886373;
publickey_row[3302] = `CIPHERTEXT_WIDTH'd5364820;
publickey_row[3303] = `CIPHERTEXT_WIDTH'd7861112;
publickey_row[3304] = `CIPHERTEXT_WIDTH'd10391910;
publickey_row[3305] = `CIPHERTEXT_WIDTH'd14595836;
publickey_row[3306] = `CIPHERTEXT_WIDTH'd13165521;
publickey_row[3307] = `CIPHERTEXT_WIDTH'd7227310;
publickey_row[3308] = `CIPHERTEXT_WIDTH'd15799618;
publickey_row[3309] = `CIPHERTEXT_WIDTH'd14064611;
publickey_row[3310] = `CIPHERTEXT_WIDTH'd11428450;
publickey_row[3311] = `CIPHERTEXT_WIDTH'd13164060;
publickey_row[3312] = `CIPHERTEXT_WIDTH'd1233503;
publickey_row[3313] = `CIPHERTEXT_WIDTH'd9053721;
publickey_row[3314] = `CIPHERTEXT_WIDTH'd14463645;
publickey_row[3315] = `CIPHERTEXT_WIDTH'd13494897;
publickey_row[3316] = `CIPHERTEXT_WIDTH'd14691422;
publickey_row[3317] = `CIPHERTEXT_WIDTH'd1745197;
publickey_row[3318] = `CIPHERTEXT_WIDTH'd7399477;
publickey_row[3319] = `CIPHERTEXT_WIDTH'd11255147;
publickey_row[3320] = `CIPHERTEXT_WIDTH'd2058425;
publickey_row[3321] = `CIPHERTEXT_WIDTH'd9058836;
publickey_row[3322] = `CIPHERTEXT_WIDTH'd6407738;
publickey_row[3323] = `CIPHERTEXT_WIDTH'd13136482;
publickey_row[3324] = `CIPHERTEXT_WIDTH'd15978509;
publickey_row[3325] = `CIPHERTEXT_WIDTH'd12228785;
publickey_row[3326] = `CIPHERTEXT_WIDTH'd14188436;
publickey_row[3327] = `CIPHERTEXT_WIDTH'd4825677;
publickey_row[3328] = `CIPHERTEXT_WIDTH'd7116302;
publickey_row[3329] = `CIPHERTEXT_WIDTH'd3172896;
publickey_row[3330] = `CIPHERTEXT_WIDTH'd3192174;
publickey_row[3331] = `CIPHERTEXT_WIDTH'd7264018;
publickey_row[3332] = `CIPHERTEXT_WIDTH'd15253428;
publickey_row[3333] = `CIPHERTEXT_WIDTH'd7208427;
publickey_row[3334] = `CIPHERTEXT_WIDTH'd11388752;
publickey_row[3335] = `CIPHERTEXT_WIDTH'd3670966;
publickey_row[3336] = `CIPHERTEXT_WIDTH'd4847737;
publickey_row[3337] = `CIPHERTEXT_WIDTH'd4322056;
publickey_row[3338] = `CIPHERTEXT_WIDTH'd8142966;
publickey_row[3339] = `CIPHERTEXT_WIDTH'd3552051;
publickey_row[3340] = `CIPHERTEXT_WIDTH'd11375547;
publickey_row[3341] = `CIPHERTEXT_WIDTH'd16681232;
publickey_row[3342] = `CIPHERTEXT_WIDTH'd13790952;
publickey_row[3343] = `CIPHERTEXT_WIDTH'd10688890;
publickey_row[3344] = `CIPHERTEXT_WIDTH'd16555785;
publickey_row[3345] = `CIPHERTEXT_WIDTH'd6899707;
publickey_row[3346] = `CIPHERTEXT_WIDTH'd15477656;
publickey_row[3347] = `CIPHERTEXT_WIDTH'd5130486;
publickey_row[3348] = `CIPHERTEXT_WIDTH'd6908757;
publickey_row[3349] = `CIPHERTEXT_WIDTH'd15614566;
publickey_row[3350] = `CIPHERTEXT_WIDTH'd7917811;
publickey_row[3351] = `CIPHERTEXT_WIDTH'd4151645;
publickey_row[3352] = `CIPHERTEXT_WIDTH'd2311046;
publickey_row[3353] = `CIPHERTEXT_WIDTH'd265322;
publickey_row[3354] = `CIPHERTEXT_WIDTH'd605218;
publickey_row[3355] = `CIPHERTEXT_WIDTH'd10348291;
publickey_row[3356] = `CIPHERTEXT_WIDTH'd12886415;
publickey_row[3357] = `CIPHERTEXT_WIDTH'd4854577;
publickey_row[3358] = `CIPHERTEXT_WIDTH'd2321067;
publickey_row[3359] = `CIPHERTEXT_WIDTH'd6018411;
publickey_row[3360] = `CIPHERTEXT_WIDTH'd4581673;
publickey_row[3361] = `CIPHERTEXT_WIDTH'd13683508;
publickey_row[3362] = `CIPHERTEXT_WIDTH'd3530071;
publickey_row[3363] = `CIPHERTEXT_WIDTH'd2746321;
publickey_row[3364] = `CIPHERTEXT_WIDTH'd7928025;
publickey_row[3365] = `CIPHERTEXT_WIDTH'd1032253;
publickey_row[3366] = `CIPHERTEXT_WIDTH'd12112111;
publickey_row[3367] = `CIPHERTEXT_WIDTH'd371527;
publickey_row[3368] = `CIPHERTEXT_WIDTH'd15558417;
publickey_row[3369] = `CIPHERTEXT_WIDTH'd10176486;
publickey_row[3370] = `CIPHERTEXT_WIDTH'd14302046;
publickey_row[3371] = `CIPHERTEXT_WIDTH'd15715632;
publickey_row[3372] = `CIPHERTEXT_WIDTH'd15384449;
publickey_row[3373] = `CIPHERTEXT_WIDTH'd5581402;
publickey_row[3374] = `CIPHERTEXT_WIDTH'd8076837;
publickey_row[3375] = `CIPHERTEXT_WIDTH'd16041852;
publickey_row[3376] = `CIPHERTEXT_WIDTH'd1544030;
publickey_row[3377] = `CIPHERTEXT_WIDTH'd11007098;
publickey_row[3378] = `CIPHERTEXT_WIDTH'd8746287;
publickey_row[3379] = `CIPHERTEXT_WIDTH'd6514091;
publickey_row[3380] = `CIPHERTEXT_WIDTH'd10793202;
publickey_row[3381] = `CIPHERTEXT_WIDTH'd14276080;
publickey_row[3382] = `CIPHERTEXT_WIDTH'd13385761;
publickey_row[3383] = `CIPHERTEXT_WIDTH'd11288475;
publickey_row[3384] = `CIPHERTEXT_WIDTH'd4957165;
publickey_row[3385] = `CIPHERTEXT_WIDTH'd11247895;
publickey_row[3386] = `CIPHERTEXT_WIDTH'd4266312;
publickey_row[3387] = `CIPHERTEXT_WIDTH'd2838100;
publickey_row[3388] = `CIPHERTEXT_WIDTH'd7552983;
publickey_row[3389] = `CIPHERTEXT_WIDTH'd14464562;
publickey_row[3390] = `CIPHERTEXT_WIDTH'd15485046;
publickey_row[3391] = `CIPHERTEXT_WIDTH'd2225410;
publickey_row[3392] = `CIPHERTEXT_WIDTH'd5265534;
publickey_row[3393] = `CIPHERTEXT_WIDTH'd3445998;
publickey_row[3394] = `CIPHERTEXT_WIDTH'd319869;
publickey_row[3395] = `CIPHERTEXT_WIDTH'd15545383;
publickey_row[3396] = `CIPHERTEXT_WIDTH'd4952812;
publickey_row[3397] = `CIPHERTEXT_WIDTH'd16327988;
publickey_row[3398] = `CIPHERTEXT_WIDTH'd10015166;
publickey_row[3399] = `CIPHERTEXT_WIDTH'd14658620;
publickey_row[3400] = `CIPHERTEXT_WIDTH'd410698;
publickey_row[3401] = `CIPHERTEXT_WIDTH'd5123037;
publickey_row[3402] = `CIPHERTEXT_WIDTH'd14272552;
publickey_row[3403] = `CIPHERTEXT_WIDTH'd15541160;
publickey_row[3404] = `CIPHERTEXT_WIDTH'd6582750;
publickey_row[3405] = `CIPHERTEXT_WIDTH'd10491702;
publickey_row[3406] = `CIPHERTEXT_WIDTH'd9938521;
publickey_row[3407] = `CIPHERTEXT_WIDTH'd11464035;
publickey_row[3408] = `CIPHERTEXT_WIDTH'd15204241;
publickey_row[3409] = `CIPHERTEXT_WIDTH'd9828753;
publickey_row[3410] = `CIPHERTEXT_WIDTH'd14266163;
publickey_row[3411] = `CIPHERTEXT_WIDTH'd13012781;
publickey_row[3412] = `CIPHERTEXT_WIDTH'd14753346;
publickey_row[3413] = `CIPHERTEXT_WIDTH'd5681115;
publickey_row[3414] = `CIPHERTEXT_WIDTH'd3109492;
publickey_row[3415] = `CIPHERTEXT_WIDTH'd4442402;
publickey_row[3416] = `CIPHERTEXT_WIDTH'd4251292;
publickey_row[3417] = `CIPHERTEXT_WIDTH'd3636371;
publickey_row[3418] = `CIPHERTEXT_WIDTH'd12528471;
publickey_row[3419] = `CIPHERTEXT_WIDTH'd15514487;
publickey_row[3420] = `CIPHERTEXT_WIDTH'd3057324;
publickey_row[3421] = `CIPHERTEXT_WIDTH'd58092;
publickey_row[3422] = `CIPHERTEXT_WIDTH'd15040169;
publickey_row[3423] = `CIPHERTEXT_WIDTH'd9582447;
publickey_row[3424] = `CIPHERTEXT_WIDTH'd13011451;
publickey_row[3425] = `CIPHERTEXT_WIDTH'd9762075;
publickey_row[3426] = `CIPHERTEXT_WIDTH'd11212733;
publickey_row[3427] = `CIPHERTEXT_WIDTH'd13922063;
publickey_row[3428] = `CIPHERTEXT_WIDTH'd1578057;
publickey_row[3429] = `CIPHERTEXT_WIDTH'd8355181;
publickey_row[3430] = `CIPHERTEXT_WIDTH'd6935502;
publickey_row[3431] = `CIPHERTEXT_WIDTH'd11293930;
publickey_row[3432] = `CIPHERTEXT_WIDTH'd13160768;
publickey_row[3433] = `CIPHERTEXT_WIDTH'd11555637;
publickey_row[3434] = `CIPHERTEXT_WIDTH'd15614386;
publickey_row[3435] = `CIPHERTEXT_WIDTH'd10521803;
publickey_row[3436] = `CIPHERTEXT_WIDTH'd13709652;
publickey_row[3437] = `CIPHERTEXT_WIDTH'd15008607;
publickey_row[3438] = `CIPHERTEXT_WIDTH'd3715790;
publickey_row[3439] = `CIPHERTEXT_WIDTH'd2075715;
publickey_row[3440] = `CIPHERTEXT_WIDTH'd16484585;
publickey_row[3441] = `CIPHERTEXT_WIDTH'd7334653;
publickey_row[3442] = `CIPHERTEXT_WIDTH'd997768;
publickey_row[3443] = `CIPHERTEXT_WIDTH'd14053143;
publickey_row[3444] = `CIPHERTEXT_WIDTH'd15956519;
publickey_row[3445] = `CIPHERTEXT_WIDTH'd14452048;
publickey_row[3446] = `CIPHERTEXT_WIDTH'd2379553;
publickey_row[3447] = `CIPHERTEXT_WIDTH'd15309203;
publickey_row[3448] = `CIPHERTEXT_WIDTH'd4613528;
publickey_row[3449] = `CIPHERTEXT_WIDTH'd5014310;
publickey_row[3450] = `CIPHERTEXT_WIDTH'd16741039;
publickey_row[3451] = `CIPHERTEXT_WIDTH'd10533053;
publickey_row[3452] = `CIPHERTEXT_WIDTH'd802552;
publickey_row[3453] = `CIPHERTEXT_WIDTH'd5848214;
publickey_row[3454] = `CIPHERTEXT_WIDTH'd11462321;
publickey_row[3455] = `CIPHERTEXT_WIDTH'd6161067;
publickey_row[3456] = `CIPHERTEXT_WIDTH'd9711128;
publickey_row[3457] = `CIPHERTEXT_WIDTH'd15431927;
publickey_row[3458] = `CIPHERTEXT_WIDTH'd4500398;
publickey_row[3459] = `CIPHERTEXT_WIDTH'd16001519;
publickey_row[3460] = `CIPHERTEXT_WIDTH'd9647160;
publickey_row[3461] = `CIPHERTEXT_WIDTH'd765252;
publickey_row[3462] = `CIPHERTEXT_WIDTH'd3876770;
publickey_row[3463] = `CIPHERTEXT_WIDTH'd15789783;
publickey_row[3464] = `CIPHERTEXT_WIDTH'd9259863;
publickey_row[3465] = `CIPHERTEXT_WIDTH'd10117952;
publickey_row[3466] = `CIPHERTEXT_WIDTH'd1979142;
publickey_row[3467] = `CIPHERTEXT_WIDTH'd6347434;
publickey_row[3468] = `CIPHERTEXT_WIDTH'd5335633;
publickey_row[3469] = `CIPHERTEXT_WIDTH'd15096426;
publickey_row[3470] = `CIPHERTEXT_WIDTH'd5867604;
publickey_row[3471] = `CIPHERTEXT_WIDTH'd14124682;
publickey_row[3472] = `CIPHERTEXT_WIDTH'd5804638;
publickey_row[3473] = `CIPHERTEXT_WIDTH'd7420522;
publickey_row[3474] = `CIPHERTEXT_WIDTH'd16606207;
publickey_row[3475] = `CIPHERTEXT_WIDTH'd1596564;
publickey_row[3476] = `CIPHERTEXT_WIDTH'd15520130;
publickey_row[3477] = `CIPHERTEXT_WIDTH'd5529894;
publickey_row[3478] = `CIPHERTEXT_WIDTH'd5860341;
publickey_row[3479] = `CIPHERTEXT_WIDTH'd15325869;
publickey_row[3480] = `CIPHERTEXT_WIDTH'd7806062;
publickey_row[3481] = `CIPHERTEXT_WIDTH'd9963592;
publickey_row[3482] = `CIPHERTEXT_WIDTH'd2175800;
publickey_row[3483] = `CIPHERTEXT_WIDTH'd6913708;
publickey_row[3484] = `CIPHERTEXT_WIDTH'd12901488;
publickey_row[3485] = `CIPHERTEXT_WIDTH'd10082885;
publickey_row[3486] = `CIPHERTEXT_WIDTH'd7696240;
publickey_row[3487] = `CIPHERTEXT_WIDTH'd5562031;
publickey_row[3488] = `CIPHERTEXT_WIDTH'd15831469;
publickey_row[3489] = `CIPHERTEXT_WIDTH'd1424032;
publickey_row[3490] = `CIPHERTEXT_WIDTH'd12664877;
publickey_row[3491] = `CIPHERTEXT_WIDTH'd4143992;
publickey_row[3492] = `CIPHERTEXT_WIDTH'd340625;
publickey_row[3493] = `CIPHERTEXT_WIDTH'd15109867;
publickey_row[3494] = `CIPHERTEXT_WIDTH'd9179072;
publickey_row[3495] = `CIPHERTEXT_WIDTH'd13030044;
publickey_row[3496] = `CIPHERTEXT_WIDTH'd13494571;
publickey_row[3497] = `CIPHERTEXT_WIDTH'd9332579;
publickey_row[3498] = `CIPHERTEXT_WIDTH'd14850620;
publickey_row[3499] = `CIPHERTEXT_WIDTH'd12414862;
publickey_row[3500] = `CIPHERTEXT_WIDTH'd8774935;
publickey_row[3501] = `CIPHERTEXT_WIDTH'd11309735;
publickey_row[3502] = `CIPHERTEXT_WIDTH'd215146;
publickey_row[3503] = `CIPHERTEXT_WIDTH'd3690174;
publickey_row[3504] = `CIPHERTEXT_WIDTH'd14049221;
publickey_row[3505] = `CIPHERTEXT_WIDTH'd12682859;
publickey_row[3506] = `CIPHERTEXT_WIDTH'd11443925;
publickey_row[3507] = `CIPHERTEXT_WIDTH'd6357099;
publickey_row[3508] = `CIPHERTEXT_WIDTH'd16649042;
publickey_row[3509] = `CIPHERTEXT_WIDTH'd9740476;
publickey_row[3510] = `CIPHERTEXT_WIDTH'd7361111;
publickey_row[3511] = `CIPHERTEXT_WIDTH'd14009322;
publickey_row[3512] = `CIPHERTEXT_WIDTH'd4535622;
publickey_row[3513] = `CIPHERTEXT_WIDTH'd1760305;
publickey_row[3514] = `CIPHERTEXT_WIDTH'd2228949;
publickey_row[3515] = `CIPHERTEXT_WIDTH'd1473653;
publickey_row[3516] = `CIPHERTEXT_WIDTH'd28561;
publickey_row[3517] = `CIPHERTEXT_WIDTH'd10308286;
publickey_row[3518] = `CIPHERTEXT_WIDTH'd11889929;
publickey_row[3519] = `CIPHERTEXT_WIDTH'd14291166;
publickey_row[3520] = `CIPHERTEXT_WIDTH'd6398600;
publickey_row[3521] = `CIPHERTEXT_WIDTH'd15088020;
publickey_row[3522] = `CIPHERTEXT_WIDTH'd12684392;
publickey_row[3523] = `CIPHERTEXT_WIDTH'd5243131;
publickey_row[3524] = `CIPHERTEXT_WIDTH'd15831551;
publickey_row[3525] = `CIPHERTEXT_WIDTH'd3339754;
publickey_row[3526] = `CIPHERTEXT_WIDTH'd10771920;
publickey_row[3527] = `CIPHERTEXT_WIDTH'd2629600;
publickey_row[3528] = `CIPHERTEXT_WIDTH'd14454409;
publickey_row[3529] = `CIPHERTEXT_WIDTH'd6979958;
publickey_row[3530] = `CIPHERTEXT_WIDTH'd2987174;
publickey_row[3531] = `CIPHERTEXT_WIDTH'd16382920;
publickey_row[3532] = `CIPHERTEXT_WIDTH'd7690655;
publickey_row[3533] = `CIPHERTEXT_WIDTH'd14229508;
publickey_row[3534] = `CIPHERTEXT_WIDTH'd10358028;
publickey_row[3535] = `CIPHERTEXT_WIDTH'd10207300;
publickey_row[3536] = `CIPHERTEXT_WIDTH'd7218458;
publickey_row[3537] = `CIPHERTEXT_WIDTH'd8598313;
publickey_row[3538] = `CIPHERTEXT_WIDTH'd798445;
publickey_row[3539] = `CIPHERTEXT_WIDTH'd6692833;
publickey_row[3540] = `CIPHERTEXT_WIDTH'd1343503;
publickey_row[3541] = `CIPHERTEXT_WIDTH'd1036446;
publickey_row[3542] = `CIPHERTEXT_WIDTH'd8438614;
publickey_row[3543] = `CIPHERTEXT_WIDTH'd9686289;
publickey_row[3544] = `CIPHERTEXT_WIDTH'd13075962;
publickey_row[3545] = `CIPHERTEXT_WIDTH'd7297491;
publickey_row[3546] = `CIPHERTEXT_WIDTH'd5106735;
publickey_row[3547] = `CIPHERTEXT_WIDTH'd9226247;
publickey_row[3548] = `CIPHERTEXT_WIDTH'd8653267;
publickey_row[3549] = `CIPHERTEXT_WIDTH'd6990863;
publickey_row[3550] = `CIPHERTEXT_WIDTH'd7915217;
publickey_row[3551] = `CIPHERTEXT_WIDTH'd12380016;
publickey_row[3552] = `CIPHERTEXT_WIDTH'd1593566;
publickey_row[3553] = `CIPHERTEXT_WIDTH'd15244784;
publickey_row[3554] = `CIPHERTEXT_WIDTH'd1937531;
publickey_row[3555] = `CIPHERTEXT_WIDTH'd3881287;
publickey_row[3556] = `CIPHERTEXT_WIDTH'd3102699;
publickey_row[3557] = `CIPHERTEXT_WIDTH'd14156727;
publickey_row[3558] = `CIPHERTEXT_WIDTH'd5593142;
publickey_row[3559] = `CIPHERTEXT_WIDTH'd15831247;
publickey_row[3560] = `CIPHERTEXT_WIDTH'd11378751;
publickey_row[3561] = `CIPHERTEXT_WIDTH'd29084;
publickey_row[3562] = `CIPHERTEXT_WIDTH'd1573473;
publickey_row[3563] = `CIPHERTEXT_WIDTH'd14954710;
publickey_row[3564] = `CIPHERTEXT_WIDTH'd5093845;
publickey_row[3565] = `CIPHERTEXT_WIDTH'd1689595;
publickey_row[3566] = `CIPHERTEXT_WIDTH'd11815197;
publickey_row[3567] = `CIPHERTEXT_WIDTH'd4137636;
publickey_row[3568] = `CIPHERTEXT_WIDTH'd15967829;
publickey_row[3569] = `CIPHERTEXT_WIDTH'd16177753;
publickey_row[3570] = `CIPHERTEXT_WIDTH'd464647;
publickey_row[3571] = `CIPHERTEXT_WIDTH'd6549374;
publickey_row[3572] = `CIPHERTEXT_WIDTH'd3943939;
publickey_row[3573] = `CIPHERTEXT_WIDTH'd7216835;
publickey_row[3574] = `CIPHERTEXT_WIDTH'd13504530;
publickey_row[3575] = `CIPHERTEXT_WIDTH'd13450810;
publickey_row[3576] = `CIPHERTEXT_WIDTH'd16748218;
publickey_row[3577] = `CIPHERTEXT_WIDTH'd15729799;
publickey_row[3578] = `CIPHERTEXT_WIDTH'd11072276;
publickey_row[3579] = `CIPHERTEXT_WIDTH'd6339150;
publickey_row[3580] = `CIPHERTEXT_WIDTH'd3117086;
publickey_row[3581] = `CIPHERTEXT_WIDTH'd4768196;
publickey_row[3582] = `CIPHERTEXT_WIDTH'd7525206;
publickey_row[3583] = `CIPHERTEXT_WIDTH'd7121745;
publickey_row[3584] = `CIPHERTEXT_WIDTH'd6097003;
publickey_row[3585] = `CIPHERTEXT_WIDTH'd4672360;
publickey_row[3586] = `CIPHERTEXT_WIDTH'd13808295;
publickey_row[3587] = `CIPHERTEXT_WIDTH'd9563433;
publickey_row[3588] = `CIPHERTEXT_WIDTH'd2942816;
publickey_row[3589] = `CIPHERTEXT_WIDTH'd3181829;
publickey_row[3590] = `CIPHERTEXT_WIDTH'd6360803;
publickey_row[3591] = `CIPHERTEXT_WIDTH'd14703175;
publickey_row[3592] = `CIPHERTEXT_WIDTH'd1684147;
publickey_row[3593] = `CIPHERTEXT_WIDTH'd11578766;
publickey_row[3594] = `CIPHERTEXT_WIDTH'd5404629;
publickey_row[3595] = `CIPHERTEXT_WIDTH'd147910;
publickey_row[3596] = `CIPHERTEXT_WIDTH'd5174547;
publickey_row[3597] = `CIPHERTEXT_WIDTH'd4692208;
publickey_row[3598] = `CIPHERTEXT_WIDTH'd8668562;
publickey_row[3599] = `CIPHERTEXT_WIDTH'd10608832;
publickey_row[3600] = `CIPHERTEXT_WIDTH'd3710240;
publickey_row[3601] = `CIPHERTEXT_WIDTH'd12528360;
publickey_row[3602] = `CIPHERTEXT_WIDTH'd2202707;
publickey_row[3603] = `CIPHERTEXT_WIDTH'd15490562;
publickey_row[3604] = `CIPHERTEXT_WIDTH'd806020;
publickey_row[3605] = `CIPHERTEXT_WIDTH'd3610370;
publickey_row[3606] = `CIPHERTEXT_WIDTH'd12458467;
publickey_row[3607] = `CIPHERTEXT_WIDTH'd6910783;
publickey_row[3608] = `CIPHERTEXT_WIDTH'd5951187;
publickey_row[3609] = `CIPHERTEXT_WIDTH'd9870159;
publickey_row[3610] = `CIPHERTEXT_WIDTH'd9082032;
publickey_row[3611] = `CIPHERTEXT_WIDTH'd4529781;
publickey_row[3612] = `CIPHERTEXT_WIDTH'd2976768;
publickey_row[3613] = `CIPHERTEXT_WIDTH'd10036289;
publickey_row[3614] = `CIPHERTEXT_WIDTH'd9966819;
publickey_row[3615] = `CIPHERTEXT_WIDTH'd7483417;
publickey_row[3616] = `CIPHERTEXT_WIDTH'd13081804;
publickey_row[3617] = `CIPHERTEXT_WIDTH'd501729;
publickey_row[3618] = `CIPHERTEXT_WIDTH'd2913361;
publickey_row[3619] = `CIPHERTEXT_WIDTH'd11233993;
publickey_row[3620] = `CIPHERTEXT_WIDTH'd14524689;
publickey_row[3621] = `CIPHERTEXT_WIDTH'd14568076;
publickey_row[3622] = `CIPHERTEXT_WIDTH'd2386306;
publickey_row[3623] = `CIPHERTEXT_WIDTH'd1740032;
publickey_row[3624] = `CIPHERTEXT_WIDTH'd8413117;
publickey_row[3625] = `CIPHERTEXT_WIDTH'd606879;
publickey_row[3626] = `CIPHERTEXT_WIDTH'd3364828;
publickey_row[3627] = `CIPHERTEXT_WIDTH'd15185311;
publickey_row[3628] = `CIPHERTEXT_WIDTH'd10968738;
publickey_row[3629] = `CIPHERTEXT_WIDTH'd16451308;
publickey_row[3630] = `CIPHERTEXT_WIDTH'd12356596;
publickey_row[3631] = `CIPHERTEXT_WIDTH'd2287346;
publickey_row[3632] = `CIPHERTEXT_WIDTH'd13751962;
publickey_row[3633] = `CIPHERTEXT_WIDTH'd6932301;
publickey_row[3634] = `CIPHERTEXT_WIDTH'd13463933;
publickey_row[3635] = `CIPHERTEXT_WIDTH'd168142;
publickey_row[3636] = `CIPHERTEXT_WIDTH'd9636756;
publickey_row[3637] = `CIPHERTEXT_WIDTH'd5034976;
publickey_row[3638] = `CIPHERTEXT_WIDTH'd5841715;
publickey_row[3639] = `CIPHERTEXT_WIDTH'd10745457;
publickey_row[3640] = `CIPHERTEXT_WIDTH'd16011385;
publickey_row[3641] = `CIPHERTEXT_WIDTH'd13435544;
publickey_row[3642] = `CIPHERTEXT_WIDTH'd4111999;
publickey_row[3643] = `CIPHERTEXT_WIDTH'd14048569;
publickey_row[3644] = `CIPHERTEXT_WIDTH'd5784473;
publickey_row[3645] = `CIPHERTEXT_WIDTH'd9612888;
publickey_row[3646] = `CIPHERTEXT_WIDTH'd3874286;
publickey_row[3647] = `CIPHERTEXT_WIDTH'd13815928;
publickey_row[3648] = `CIPHERTEXT_WIDTH'd11530435;
publickey_row[3649] = `CIPHERTEXT_WIDTH'd16090161;
publickey_row[3650] = `CIPHERTEXT_WIDTH'd11160514;
publickey_row[3651] = `CIPHERTEXT_WIDTH'd14403089;
publickey_row[3652] = `CIPHERTEXT_WIDTH'd14764398;
publickey_row[3653] = `CIPHERTEXT_WIDTH'd13407552;
publickey_row[3654] = `CIPHERTEXT_WIDTH'd12814400;
publickey_row[3655] = `CIPHERTEXT_WIDTH'd8962552;
publickey_row[3656] = `CIPHERTEXT_WIDTH'd6339734;
publickey_row[3657] = `CIPHERTEXT_WIDTH'd11994754;
publickey_row[3658] = `CIPHERTEXT_WIDTH'd9072918;
publickey_row[3659] = `CIPHERTEXT_WIDTH'd16480276;
publickey_row[3660] = `CIPHERTEXT_WIDTH'd8419141;
publickey_row[3661] = `CIPHERTEXT_WIDTH'd14323763;
publickey_row[3662] = `CIPHERTEXT_WIDTH'd8488299;
publickey_row[3663] = `CIPHERTEXT_WIDTH'd3256775;
publickey_row[3664] = `CIPHERTEXT_WIDTH'd11644471;
publickey_row[3665] = `CIPHERTEXT_WIDTH'd4041362;
publickey_row[3666] = `CIPHERTEXT_WIDTH'd7480109;
publickey_row[3667] = `CIPHERTEXT_WIDTH'd7868476;
publickey_row[3668] = `CIPHERTEXT_WIDTH'd12366954;
publickey_row[3669] = `CIPHERTEXT_WIDTH'd2055277;
publickey_row[3670] = `CIPHERTEXT_WIDTH'd10863402;
publickey_row[3671] = `CIPHERTEXT_WIDTH'd3218861;
publickey_row[3672] = `CIPHERTEXT_WIDTH'd6329883;
publickey_row[3673] = `CIPHERTEXT_WIDTH'd3510959;
publickey_row[3674] = `CIPHERTEXT_WIDTH'd692687;
publickey_row[3675] = `CIPHERTEXT_WIDTH'd1822341;
publickey_row[3676] = `CIPHERTEXT_WIDTH'd10057721;
publickey_row[3677] = `CIPHERTEXT_WIDTH'd5097504;
publickey_row[3678] = `CIPHERTEXT_WIDTH'd7869713;
publickey_row[3679] = `CIPHERTEXT_WIDTH'd897344;
publickey_row[3680] = `CIPHERTEXT_WIDTH'd4899053;
publickey_row[3681] = `CIPHERTEXT_WIDTH'd3415676;
publickey_row[3682] = `CIPHERTEXT_WIDTH'd4469748;
publickey_row[3683] = `CIPHERTEXT_WIDTH'd14393200;
publickey_row[3684] = `CIPHERTEXT_WIDTH'd6676662;
publickey_row[3685] = `CIPHERTEXT_WIDTH'd8468884;
publickey_row[3686] = `CIPHERTEXT_WIDTH'd5745607;
publickey_row[3687] = `CIPHERTEXT_WIDTH'd7804754;
publickey_row[3688] = `CIPHERTEXT_WIDTH'd16090133;
publickey_row[3689] = `CIPHERTEXT_WIDTH'd13291902;
publickey_row[3690] = `CIPHERTEXT_WIDTH'd5935024;
publickey_row[3691] = `CIPHERTEXT_WIDTH'd2329983;
publickey_row[3692] = `CIPHERTEXT_WIDTH'd11630531;
publickey_row[3693] = `CIPHERTEXT_WIDTH'd14321356;
publickey_row[3694] = `CIPHERTEXT_WIDTH'd14809958;
publickey_row[3695] = `CIPHERTEXT_WIDTH'd5953186;
publickey_row[3696] = `CIPHERTEXT_WIDTH'd4746330;
publickey_row[3697] = `CIPHERTEXT_WIDTH'd4734402;
publickey_row[3698] = `CIPHERTEXT_WIDTH'd3213304;
publickey_row[3699] = `CIPHERTEXT_WIDTH'd10131140;
publickey_row[3700] = `CIPHERTEXT_WIDTH'd14759238;
publickey_row[3701] = `CIPHERTEXT_WIDTH'd853038;
publickey_row[3702] = `CIPHERTEXT_WIDTH'd1562020;
publickey_row[3703] = `CIPHERTEXT_WIDTH'd876164;
publickey_row[3704] = `CIPHERTEXT_WIDTH'd8005046;
publickey_row[3705] = `CIPHERTEXT_WIDTH'd8265590;
publickey_row[3706] = `CIPHERTEXT_WIDTH'd16215429;
publickey_row[3707] = `CIPHERTEXT_WIDTH'd9501373;
publickey_row[3708] = `CIPHERTEXT_WIDTH'd10697081;
publickey_row[3709] = `CIPHERTEXT_WIDTH'd11716272;
publickey_row[3710] = `CIPHERTEXT_WIDTH'd15797805;
publickey_row[3711] = `CIPHERTEXT_WIDTH'd9342426;
publickey_row[3712] = `CIPHERTEXT_WIDTH'd4294370;
publickey_row[3713] = `CIPHERTEXT_WIDTH'd4202443;
publickey_row[3714] = `CIPHERTEXT_WIDTH'd4905933;
publickey_row[3715] = `CIPHERTEXT_WIDTH'd897670;
publickey_row[3716] = `CIPHERTEXT_WIDTH'd5228786;
publickey_row[3717] = `CIPHERTEXT_WIDTH'd7822644;
publickey_row[3718] = `CIPHERTEXT_WIDTH'd11617312;
publickey_row[3719] = `CIPHERTEXT_WIDTH'd12633090;
publickey_row[3720] = `CIPHERTEXT_WIDTH'd3018853;
publickey_row[3721] = `CIPHERTEXT_WIDTH'd6193201;
publickey_row[3722] = `CIPHERTEXT_WIDTH'd10423798;
publickey_row[3723] = `CIPHERTEXT_WIDTH'd12550487;
publickey_row[3724] = `CIPHERTEXT_WIDTH'd11187976;
publickey_row[3725] = `CIPHERTEXT_WIDTH'd5259340;
publickey_row[3726] = `CIPHERTEXT_WIDTH'd224089;
publickey_row[3727] = `CIPHERTEXT_WIDTH'd3351653;
publickey_row[3728] = `CIPHERTEXT_WIDTH'd9193024;
publickey_row[3729] = `CIPHERTEXT_WIDTH'd5100137;
publickey_row[3730] = `CIPHERTEXT_WIDTH'd10352241;
publickey_row[3731] = `CIPHERTEXT_WIDTH'd4227108;
publickey_row[3732] = `CIPHERTEXT_WIDTH'd10696303;
publickey_row[3733] = `CIPHERTEXT_WIDTH'd6670489;
publickey_row[3734] = `CIPHERTEXT_WIDTH'd16437185;
publickey_row[3735] = `CIPHERTEXT_WIDTH'd3350376;
publickey_row[3736] = `CIPHERTEXT_WIDTH'd2910701;
publickey_row[3737] = `CIPHERTEXT_WIDTH'd8037114;
publickey_row[3738] = `CIPHERTEXT_WIDTH'd8687774;
publickey_row[3739] = `CIPHERTEXT_WIDTH'd12540714;
publickey_row[3740] = `CIPHERTEXT_WIDTH'd8637698;
publickey_row[3741] = `CIPHERTEXT_WIDTH'd540952;
publickey_row[3742] = `CIPHERTEXT_WIDTH'd14132857;
publickey_row[3743] = `CIPHERTEXT_WIDTH'd909763;
publickey_row[3744] = `CIPHERTEXT_WIDTH'd14355708;
publickey_row[3745] = `CIPHERTEXT_WIDTH'd11840400;
publickey_row[3746] = `CIPHERTEXT_WIDTH'd11449898;
publickey_row[3747] = `CIPHERTEXT_WIDTH'd11226017;
publickey_row[3748] = `CIPHERTEXT_WIDTH'd2469233;
publickey_row[3749] = `CIPHERTEXT_WIDTH'd6032571;
publickey_row[3750] = `CIPHERTEXT_WIDTH'd15838925;
publickey_row[3751] = `CIPHERTEXT_WIDTH'd9154015;
publickey_row[3752] = `CIPHERTEXT_WIDTH'd12865573;
publickey_row[3753] = `CIPHERTEXT_WIDTH'd12010370;
publickey_row[3754] = `CIPHERTEXT_WIDTH'd5144745;
publickey_row[3755] = `CIPHERTEXT_WIDTH'd3632289;
publickey_row[3756] = `CIPHERTEXT_WIDTH'd5360986;
publickey_row[3757] = `CIPHERTEXT_WIDTH'd12885149;
publickey_row[3758] = `CIPHERTEXT_WIDTH'd12387265;
publickey_row[3759] = `CIPHERTEXT_WIDTH'd8741125;
publickey_row[3760] = `CIPHERTEXT_WIDTH'd9781473;
publickey_row[3761] = `CIPHERTEXT_WIDTH'd16025808;
publickey_row[3762] = `CIPHERTEXT_WIDTH'd6153316;
publickey_row[3763] = `CIPHERTEXT_WIDTH'd4520243;
publickey_row[3764] = `CIPHERTEXT_WIDTH'd11077217;
publickey_row[3765] = `CIPHERTEXT_WIDTH'd8098205;
publickey_row[3766] = `CIPHERTEXT_WIDTH'd3757112;
publickey_row[3767] = `CIPHERTEXT_WIDTH'd12137708;
publickey_row[3768] = `CIPHERTEXT_WIDTH'd11749379;
publickey_row[3769] = `CIPHERTEXT_WIDTH'd12306131;
publickey_row[3770] = `CIPHERTEXT_WIDTH'd16405865;
publickey_row[3771] = `CIPHERTEXT_WIDTH'd5129181;
publickey_row[3772] = `CIPHERTEXT_WIDTH'd8764039;
publickey_row[3773] = `CIPHERTEXT_WIDTH'd1248891;
publickey_row[3774] = `CIPHERTEXT_WIDTH'd9412147;
publickey_row[3775] = `CIPHERTEXT_WIDTH'd1763522;
publickey_row[3776] = `CIPHERTEXT_WIDTH'd970450;
publickey_row[3777] = `CIPHERTEXT_WIDTH'd82541;
publickey_row[3778] = `CIPHERTEXT_WIDTH'd7032630;
publickey_row[3779] = `CIPHERTEXT_WIDTH'd12028375;
publickey_row[3780] = `CIPHERTEXT_WIDTH'd2707460;
publickey_row[3781] = `CIPHERTEXT_WIDTH'd16492813;
publickey_row[3782] = `CIPHERTEXT_WIDTH'd14437428;
publickey_row[3783] = `CIPHERTEXT_WIDTH'd10196396;
publickey_row[3784] = `CIPHERTEXT_WIDTH'd14119653;
publickey_row[3785] = `CIPHERTEXT_WIDTH'd2795887;
publickey_row[3786] = `CIPHERTEXT_WIDTH'd7061941;
publickey_row[3787] = `CIPHERTEXT_WIDTH'd2493737;
publickey_row[3788] = `CIPHERTEXT_WIDTH'd595397;
publickey_row[3789] = `CIPHERTEXT_WIDTH'd1610677;
publickey_row[3790] = `CIPHERTEXT_WIDTH'd9677561;
publickey_row[3791] = `CIPHERTEXT_WIDTH'd6577583;
publickey_row[3792] = `CIPHERTEXT_WIDTH'd1869423;
publickey_row[3793] = `CIPHERTEXT_WIDTH'd8737789;
publickey_row[3794] = `CIPHERTEXT_WIDTH'd16391597;
publickey_row[3795] = `CIPHERTEXT_WIDTH'd6140009;
publickey_row[3796] = `CIPHERTEXT_WIDTH'd7128560;
publickey_row[3797] = `CIPHERTEXT_WIDTH'd15476471;
publickey_row[3798] = `CIPHERTEXT_WIDTH'd3754467;
publickey_row[3799] = `CIPHERTEXT_WIDTH'd2717786;
publickey_row[3800] = `CIPHERTEXT_WIDTH'd12923472;
publickey_row[3801] = `CIPHERTEXT_WIDTH'd1479372;
publickey_row[3802] = `CIPHERTEXT_WIDTH'd559545;
publickey_row[3803] = `CIPHERTEXT_WIDTH'd14901386;
publickey_row[3804] = `CIPHERTEXT_WIDTH'd8031435;
publickey_row[3805] = `CIPHERTEXT_WIDTH'd14137234;
publickey_row[3806] = `CIPHERTEXT_WIDTH'd13681874;
publickey_row[3807] = `CIPHERTEXT_WIDTH'd1877027;
publickey_row[3808] = `CIPHERTEXT_WIDTH'd15931568;
publickey_row[3809] = `CIPHERTEXT_WIDTH'd6874722;
publickey_row[3810] = `CIPHERTEXT_WIDTH'd16682585;
publickey_row[3811] = `CIPHERTEXT_WIDTH'd1287866;
publickey_row[3812] = `CIPHERTEXT_WIDTH'd2573233;
publickey_row[3813] = `CIPHERTEXT_WIDTH'd5547320;
publickey_row[3814] = `CIPHERTEXT_WIDTH'd5812511;
publickey_row[3815] = `CIPHERTEXT_WIDTH'd3498358;
publickey_row[3816] = `CIPHERTEXT_WIDTH'd1236647;
publickey_row[3817] = `CIPHERTEXT_WIDTH'd7851415;
publickey_row[3818] = `CIPHERTEXT_WIDTH'd10076453;
publickey_row[3819] = `CIPHERTEXT_WIDTH'd15017677;
publickey_row[3820] = `CIPHERTEXT_WIDTH'd16484810;
publickey_row[3821] = `CIPHERTEXT_WIDTH'd13710074;
publickey_row[3822] = `CIPHERTEXT_WIDTH'd2203636;
publickey_row[3823] = `CIPHERTEXT_WIDTH'd657132;
publickey_row[3824] = `CIPHERTEXT_WIDTH'd13072996;
publickey_row[3825] = `CIPHERTEXT_WIDTH'd1168319;
publickey_row[3826] = `CIPHERTEXT_WIDTH'd14588655;
publickey_row[3827] = `CIPHERTEXT_WIDTH'd5833069;
publickey_row[3828] = `CIPHERTEXT_WIDTH'd15546628;
publickey_row[3829] = `CIPHERTEXT_WIDTH'd7191008;
publickey_row[3830] = `CIPHERTEXT_WIDTH'd12422307;
publickey_row[3831] = `CIPHERTEXT_WIDTH'd16558967;
publickey_row[3832] = `CIPHERTEXT_WIDTH'd7640358;
publickey_row[3833] = `CIPHERTEXT_WIDTH'd6659783;
publickey_row[3834] = `CIPHERTEXT_WIDTH'd13440916;
publickey_row[3835] = `CIPHERTEXT_WIDTH'd8924425;
publickey_row[3836] = `CIPHERTEXT_WIDTH'd2793442;
publickey_row[3837] = `CIPHERTEXT_WIDTH'd9783224;
publickey_row[3838] = `CIPHERTEXT_WIDTH'd7968907;
publickey_row[3839] = `CIPHERTEXT_WIDTH'd10213901;
publickey_row[3840] = `CIPHERTEXT_WIDTH'd4087787;
publickey_row[3841] = `CIPHERTEXT_WIDTH'd7735064;
publickey_row[3842] = `CIPHERTEXT_WIDTH'd13621560;
publickey_row[3843] = `CIPHERTEXT_WIDTH'd3621364;
publickey_row[3844] = `CIPHERTEXT_WIDTH'd5264859;
publickey_row[3845] = `CIPHERTEXT_WIDTH'd5732067;
publickey_row[3846] = `CIPHERTEXT_WIDTH'd4385180;
publickey_row[3847] = `CIPHERTEXT_WIDTH'd12250417;
publickey_row[3848] = `CIPHERTEXT_WIDTH'd16471439;
publickey_row[3849] = `CIPHERTEXT_WIDTH'd13687237;
publickey_row[3850] = `CIPHERTEXT_WIDTH'd11018523;
publickey_row[3851] = `CIPHERTEXT_WIDTH'd5232503;
publickey_row[3852] = `CIPHERTEXT_WIDTH'd763095;
publickey_row[3853] = `CIPHERTEXT_WIDTH'd10816816;
publickey_row[3854] = `CIPHERTEXT_WIDTH'd2275646;
publickey_row[3855] = `CIPHERTEXT_WIDTH'd4484619;
publickey_row[3856] = `CIPHERTEXT_WIDTH'd11851121;
publickey_row[3857] = `CIPHERTEXT_WIDTH'd9304252;
publickey_row[3858] = `CIPHERTEXT_WIDTH'd13581777;
publickey_row[3859] = `CIPHERTEXT_WIDTH'd14055812;
publickey_row[3860] = `CIPHERTEXT_WIDTH'd9912346;
publickey_row[3861] = `CIPHERTEXT_WIDTH'd7430207;
publickey_row[3862] = `CIPHERTEXT_WIDTH'd2062638;
publickey_row[3863] = `CIPHERTEXT_WIDTH'd14261904;
publickey_row[3864] = `CIPHERTEXT_WIDTH'd3764032;
publickey_row[3865] = `CIPHERTEXT_WIDTH'd11032343;
publickey_row[3866] = `CIPHERTEXT_WIDTH'd5663242;
publickey_row[3867] = `CIPHERTEXT_WIDTH'd6233114;
publickey_row[3868] = `CIPHERTEXT_WIDTH'd3331467;
publickey_row[3869] = `CIPHERTEXT_WIDTH'd7182846;
publickey_row[3870] = `CIPHERTEXT_WIDTH'd4940047;
publickey_row[3871] = `CIPHERTEXT_WIDTH'd10043856;
publickey_row[3872] = `CIPHERTEXT_WIDTH'd3257133;
publickey_row[3873] = `CIPHERTEXT_WIDTH'd1586349;
publickey_row[3874] = `CIPHERTEXT_WIDTH'd12069289;
publickey_row[3875] = `CIPHERTEXT_WIDTH'd9785897;
publickey_row[3876] = `CIPHERTEXT_WIDTH'd6427944;
publickey_row[3877] = `CIPHERTEXT_WIDTH'd4533231;
publickey_row[3878] = `CIPHERTEXT_WIDTH'd14714434;
publickey_row[3879] = `CIPHERTEXT_WIDTH'd7901312;
publickey_row[3880] = `CIPHERTEXT_WIDTH'd13968530;
publickey_row[3881] = `CIPHERTEXT_WIDTH'd14745186;
publickey_row[3882] = `CIPHERTEXT_WIDTH'd676193;
publickey_row[3883] = `CIPHERTEXT_WIDTH'd5538117;
publickey_row[3884] = `CIPHERTEXT_WIDTH'd8925507;
publickey_row[3885] = `CIPHERTEXT_WIDTH'd5067077;
publickey_row[3886] = `CIPHERTEXT_WIDTH'd14439160;
publickey_row[3887] = `CIPHERTEXT_WIDTH'd13618179;
publickey_row[3888] = `CIPHERTEXT_WIDTH'd12757304;
publickey_row[3889] = `CIPHERTEXT_WIDTH'd11342873;
publickey_row[3890] = `CIPHERTEXT_WIDTH'd59030;
publickey_row[3891] = `CIPHERTEXT_WIDTH'd8981561;
publickey_row[3892] = `CIPHERTEXT_WIDTH'd13234455;
publickey_row[3893] = `CIPHERTEXT_WIDTH'd3398788;
publickey_row[3894] = `CIPHERTEXT_WIDTH'd15420380;
publickey_row[3895] = `CIPHERTEXT_WIDTH'd15856921;
publickey_row[3896] = `CIPHERTEXT_WIDTH'd2073919;
publickey_row[3897] = `CIPHERTEXT_WIDTH'd7404765;
publickey_row[3898] = `CIPHERTEXT_WIDTH'd14772731;
publickey_row[3899] = `CIPHERTEXT_WIDTH'd13250442;
publickey_row[3900] = `CIPHERTEXT_WIDTH'd8783761;
publickey_row[3901] = `CIPHERTEXT_WIDTH'd1696687;
publickey_row[3902] = `CIPHERTEXT_WIDTH'd10869761;
publickey_row[3903] = `CIPHERTEXT_WIDTH'd16093863;
publickey_row[3904] = `CIPHERTEXT_WIDTH'd15975933;
publickey_row[3905] = `CIPHERTEXT_WIDTH'd5781450;
publickey_row[3906] = `CIPHERTEXT_WIDTH'd15062807;
publickey_row[3907] = `CIPHERTEXT_WIDTH'd14482338;
publickey_row[3908] = `CIPHERTEXT_WIDTH'd5622818;
publickey_row[3909] = `CIPHERTEXT_WIDTH'd4364351;
publickey_row[3910] = `CIPHERTEXT_WIDTH'd10551087;
publickey_row[3911] = `CIPHERTEXT_WIDTH'd11014449;
publickey_row[3912] = `CIPHERTEXT_WIDTH'd9179586;
publickey_row[3913] = `CIPHERTEXT_WIDTH'd13929918;
publickey_row[3914] = `CIPHERTEXT_WIDTH'd2278691;
publickey_row[3915] = `CIPHERTEXT_WIDTH'd16398942;
publickey_row[3916] = `CIPHERTEXT_WIDTH'd423625;
publickey_row[3917] = `CIPHERTEXT_WIDTH'd671278;
publickey_row[3918] = `CIPHERTEXT_WIDTH'd4888546;
publickey_row[3919] = `CIPHERTEXT_WIDTH'd14604624;
publickey_row[3920] = `CIPHERTEXT_WIDTH'd1126216;
publickey_row[3921] = `CIPHERTEXT_WIDTH'd12496185;
publickey_row[3922] = `CIPHERTEXT_WIDTH'd14866623;
publickey_row[3923] = `CIPHERTEXT_WIDTH'd9951252;
publickey_row[3924] = `CIPHERTEXT_WIDTH'd3192022;
publickey_row[3925] = `CIPHERTEXT_WIDTH'd9773174;
publickey_row[3926] = `CIPHERTEXT_WIDTH'd15806073;
publickey_row[3927] = `CIPHERTEXT_WIDTH'd15766135;
publickey_row[3928] = `CIPHERTEXT_WIDTH'd2370188;
publickey_row[3929] = `CIPHERTEXT_WIDTH'd14887053;
publickey_row[3930] = `CIPHERTEXT_WIDTH'd7776339;
publickey_row[3931] = `CIPHERTEXT_WIDTH'd9769130;
publickey_row[3932] = `CIPHERTEXT_WIDTH'd2055094;
publickey_row[3933] = `CIPHERTEXT_WIDTH'd9316351;
publickey_row[3934] = `CIPHERTEXT_WIDTH'd12898830;
publickey_row[3935] = `CIPHERTEXT_WIDTH'd8079999;
publickey_row[3936] = `CIPHERTEXT_WIDTH'd1326098;
publickey_row[3937] = `CIPHERTEXT_WIDTH'd8343280;
publickey_row[3938] = `CIPHERTEXT_WIDTH'd588084;
publickey_row[3939] = `CIPHERTEXT_WIDTH'd12345429;
publickey_row[3940] = `CIPHERTEXT_WIDTH'd2210545;
publickey_row[3941] = `CIPHERTEXT_WIDTH'd1613657;
publickey_row[3942] = `CIPHERTEXT_WIDTH'd11801;
publickey_row[3943] = `CIPHERTEXT_WIDTH'd8793363;
publickey_row[3944] = `CIPHERTEXT_WIDTH'd7462032;
publickey_row[3945] = `CIPHERTEXT_WIDTH'd306829;
publickey_row[3946] = `CIPHERTEXT_WIDTH'd13534085;
publickey_row[3947] = `CIPHERTEXT_WIDTH'd8378914;
publickey_row[3948] = `CIPHERTEXT_WIDTH'd4521159;
publickey_row[3949] = `CIPHERTEXT_WIDTH'd6638002;
publickey_row[3950] = `CIPHERTEXT_WIDTH'd1465879;
publickey_row[3951] = `CIPHERTEXT_WIDTH'd4234300;
publickey_row[3952] = `CIPHERTEXT_WIDTH'd7391108;
publickey_row[3953] = `CIPHERTEXT_WIDTH'd16561671;
publickey_row[3954] = `CIPHERTEXT_WIDTH'd9974494;
publickey_row[3955] = `CIPHERTEXT_WIDTH'd1961784;
publickey_row[3956] = `CIPHERTEXT_WIDTH'd9669579;
publickey_row[3957] = `CIPHERTEXT_WIDTH'd6203866;
publickey_row[3958] = `CIPHERTEXT_WIDTH'd11927267;
publickey_row[3959] = `CIPHERTEXT_WIDTH'd15694766;
publickey_row[3960] = `CIPHERTEXT_WIDTH'd5459020;
publickey_row[3961] = `CIPHERTEXT_WIDTH'd9993138;
publickey_row[3962] = `CIPHERTEXT_WIDTH'd9141515;
publickey_row[3963] = `CIPHERTEXT_WIDTH'd2320456;
publickey_row[3964] = `CIPHERTEXT_WIDTH'd1801558;
publickey_row[3965] = `CIPHERTEXT_WIDTH'd4623858;
publickey_row[3966] = `CIPHERTEXT_WIDTH'd4506947;
publickey_row[3967] = `CIPHERTEXT_WIDTH'd1980388;
publickey_row[3968] = `CIPHERTEXT_WIDTH'd4112638;
publickey_row[3969] = `CIPHERTEXT_WIDTH'd6725117;
publickey_row[3970] = `CIPHERTEXT_WIDTH'd10376396;
publickey_row[3971] = `CIPHERTEXT_WIDTH'd569308;
publickey_row[3972] = `CIPHERTEXT_WIDTH'd7051757;
publickey_row[3973] = `CIPHERTEXT_WIDTH'd9060050;
publickey_row[3974] = `CIPHERTEXT_WIDTH'd15881436;
publickey_row[3975] = `CIPHERTEXT_WIDTH'd3098560;
publickey_row[3976] = `CIPHERTEXT_WIDTH'd16565215;
publickey_row[3977] = `CIPHERTEXT_WIDTH'd8177503;
publickey_row[3978] = `CIPHERTEXT_WIDTH'd11407828;
publickey_row[3979] = `CIPHERTEXT_WIDTH'd2962994;
publickey_row[3980] = `CIPHERTEXT_WIDTH'd16298499;
publickey_row[3981] = `CIPHERTEXT_WIDTH'd14092205;
publickey_row[3982] = `CIPHERTEXT_WIDTH'd4376054;
publickey_row[3983] = `CIPHERTEXT_WIDTH'd14800803;
publickey_row[3984] = `CIPHERTEXT_WIDTH'd2977956;
publickey_row[3985] = `CIPHERTEXT_WIDTH'd10992189;
publickey_row[3986] = `CIPHERTEXT_WIDTH'd15704020;
publickey_row[3987] = `CIPHERTEXT_WIDTH'd772878;
publickey_row[3988] = `CIPHERTEXT_WIDTH'd2753694;
publickey_row[3989] = `CIPHERTEXT_WIDTH'd10414447;
publickey_row[3990] = `CIPHERTEXT_WIDTH'd7747381;
publickey_row[3991] = `CIPHERTEXT_WIDTH'd10040771;
publickey_row[3992] = `CIPHERTEXT_WIDTH'd15109865;
publickey_row[3993] = `CIPHERTEXT_WIDTH'd2241244;
publickey_row[3994] = `CIPHERTEXT_WIDTH'd11957745;
publickey_row[3995] = `CIPHERTEXT_WIDTH'd16427843;
publickey_row[3996] = `CIPHERTEXT_WIDTH'd2560849;
publickey_row[3997] = `CIPHERTEXT_WIDTH'd7074344;
publickey_row[3998] = `CIPHERTEXT_WIDTH'd293191;
publickey_row[3999] = `CIPHERTEXT_WIDTH'd6733841;
publickey_row[4000] = `CIPHERTEXT_WIDTH'd9185119;
publickey_row[4001] = `CIPHERTEXT_WIDTH'd9055318;
publickey_row[4002] = `CIPHERTEXT_WIDTH'd12204097;
publickey_row[4003] = `CIPHERTEXT_WIDTH'd6179446;
publickey_row[4004] = `CIPHERTEXT_WIDTH'd1763138;
publickey_row[4005] = `CIPHERTEXT_WIDTH'd15767429;
publickey_row[4006] = `CIPHERTEXT_WIDTH'd4148189;
publickey_row[4007] = `CIPHERTEXT_WIDTH'd2383133;
publickey_row[4008] = `CIPHERTEXT_WIDTH'd1678527;
publickey_row[4009] = `CIPHERTEXT_WIDTH'd15975700;
publickey_row[4010] = `CIPHERTEXT_WIDTH'd8290983;
publickey_row[4011] = `CIPHERTEXT_WIDTH'd2302005;
publickey_row[4012] = `CIPHERTEXT_WIDTH'd7060621;
publickey_row[4013] = `CIPHERTEXT_WIDTH'd3817218;
publickey_row[4014] = `CIPHERTEXT_WIDTH'd7788951;
publickey_row[4015] = `CIPHERTEXT_WIDTH'd12193493;
publickey_row[4016] = `CIPHERTEXT_WIDTH'd2120436;
publickey_row[4017] = `CIPHERTEXT_WIDTH'd12062068;
publickey_row[4018] = `CIPHERTEXT_WIDTH'd9608601;
publickey_row[4019] = `CIPHERTEXT_WIDTH'd4088842;
publickey_row[4020] = `CIPHERTEXT_WIDTH'd3888212;
publickey_row[4021] = `CIPHERTEXT_WIDTH'd4154905;
publickey_row[4022] = `CIPHERTEXT_WIDTH'd6910922;
publickey_row[4023] = `CIPHERTEXT_WIDTH'd15582117;
publickey_row[4024] = `CIPHERTEXT_WIDTH'd1960643;
publickey_row[4025] = `CIPHERTEXT_WIDTH'd16395157;
publickey_row[4026] = `CIPHERTEXT_WIDTH'd14817978;
publickey_row[4027] = `CIPHERTEXT_WIDTH'd8896736;
publickey_row[4028] = `CIPHERTEXT_WIDTH'd9604594;
publickey_row[4029] = `CIPHERTEXT_WIDTH'd11034300;
publickey_row[4030] = `CIPHERTEXT_WIDTH'd9903580;
publickey_row[4031] = `CIPHERTEXT_WIDTH'd10220814;
publickey_row[4032] = `CIPHERTEXT_WIDTH'd13158897;
publickey_row[4033] = `CIPHERTEXT_WIDTH'd11513419;
publickey_row[4034] = `CIPHERTEXT_WIDTH'd3419436;
publickey_row[4035] = `CIPHERTEXT_WIDTH'd11987246;
publickey_row[4036] = `CIPHERTEXT_WIDTH'd15817218;
publickey_row[4037] = `CIPHERTEXT_WIDTH'd12284063;
publickey_row[4038] = `CIPHERTEXT_WIDTH'd6574083;
publickey_row[4039] = `CIPHERTEXT_WIDTH'd6527843;
publickey_row[4040] = `CIPHERTEXT_WIDTH'd8058076;
publickey_row[4041] = `CIPHERTEXT_WIDTH'd13384517;
publickey_row[4042] = `CIPHERTEXT_WIDTH'd13849917;
publickey_row[4043] = `CIPHERTEXT_WIDTH'd14710387;
publickey_row[4044] = `CIPHERTEXT_WIDTH'd193722;
publickey_row[4045] = `CIPHERTEXT_WIDTH'd10963032;
publickey_row[4046] = `CIPHERTEXT_WIDTH'd9982221;
publickey_row[4047] = `CIPHERTEXT_WIDTH'd15766551;
publickey_row[4048] = `CIPHERTEXT_WIDTH'd5186693;
publickey_row[4049] = `CIPHERTEXT_WIDTH'd4192728;
publickey_row[4050] = `CIPHERTEXT_WIDTH'd9750463;
publickey_row[4051] = `CIPHERTEXT_WIDTH'd10583427;
publickey_row[4052] = `CIPHERTEXT_WIDTH'd5607698;
publickey_row[4053] = `CIPHERTEXT_WIDTH'd14470823;
publickey_row[4054] = `CIPHERTEXT_WIDTH'd9831992;
publickey_row[4055] = `CIPHERTEXT_WIDTH'd6487781;
publickey_row[4056] = `CIPHERTEXT_WIDTH'd7170209;
publickey_row[4057] = `CIPHERTEXT_WIDTH'd11703679;
publickey_row[4058] = `CIPHERTEXT_WIDTH'd15971700;
publickey_row[4059] = `CIPHERTEXT_WIDTH'd9096617;
publickey_row[4060] = `CIPHERTEXT_WIDTH'd3685801;
publickey_row[4061] = `CIPHERTEXT_WIDTH'd8726368;
publickey_row[4062] = `CIPHERTEXT_WIDTH'd6379613;
publickey_row[4063] = `CIPHERTEXT_WIDTH'd3317040;
publickey_row[4064] = `CIPHERTEXT_WIDTH'd1086267;
publickey_row[4065] = `CIPHERTEXT_WIDTH'd16182007;
publickey_row[4066] = `CIPHERTEXT_WIDTH'd1897196;
publickey_row[4067] = `CIPHERTEXT_WIDTH'd13261491;
publickey_row[4068] = `CIPHERTEXT_WIDTH'd6527252;
publickey_row[4069] = `CIPHERTEXT_WIDTH'd4643231;
publickey_row[4070] = `CIPHERTEXT_WIDTH'd10749213;
publickey_row[4071] = `CIPHERTEXT_WIDTH'd6649945;
publickey_row[4072] = `CIPHERTEXT_WIDTH'd13521642;
publickey_row[4073] = `CIPHERTEXT_WIDTH'd1198952;
publickey_row[4074] = `CIPHERTEXT_WIDTH'd8835164;
publickey_row[4075] = `CIPHERTEXT_WIDTH'd14018172;
publickey_row[4076] = `CIPHERTEXT_WIDTH'd3549435;
publickey_row[4077] = `CIPHERTEXT_WIDTH'd2190272;
publickey_row[4078] = `CIPHERTEXT_WIDTH'd12309539;
publickey_row[4079] = `CIPHERTEXT_WIDTH'd8229472;
publickey_row[4080] = `CIPHERTEXT_WIDTH'd13781123;
publickey_row[4081] = `CIPHERTEXT_WIDTH'd561684;
publickey_row[4082] = `CIPHERTEXT_WIDTH'd9797635;
publickey_row[4083] = `CIPHERTEXT_WIDTH'd4026885;
publickey_row[4084] = `CIPHERTEXT_WIDTH'd7425015;
publickey_row[4085] = `CIPHERTEXT_WIDTH'd9807580;
publickey_row[4086] = `CIPHERTEXT_WIDTH'd13777379;
publickey_row[4087] = `CIPHERTEXT_WIDTH'd13125432;
publickey_row[4088] = `CIPHERTEXT_WIDTH'd15856717;
publickey_row[4089] = `CIPHERTEXT_WIDTH'd9815702;
publickey_row[4090] = `CIPHERTEXT_WIDTH'd16212141;
publickey_row[4091] = `CIPHERTEXT_WIDTH'd10634932;
publickey_row[4092] = `CIPHERTEXT_WIDTH'd9334235;
publickey_row[4093] = `CIPHERTEXT_WIDTH'd4713793;
publickey_row[4094] = `CIPHERTEXT_WIDTH'd13377975;
publickey_row[4095] = `CIPHERTEXT_WIDTH'd3675263;
publickey_row[4096] = `CIPHERTEXT_WIDTH'd14890871;
publickey_row[4097] = `CIPHERTEXT_WIDTH'd8156437;
publickey_row[4098] = `CIPHERTEXT_WIDTH'd11207240;
publickey_row[4099] = `CIPHERTEXT_WIDTH'd350790;
publickey_row[4100] = `CIPHERTEXT_WIDTH'd3681415;
publickey_row[4101] = `CIPHERTEXT_WIDTH'd4291413;
publickey_row[4102] = `CIPHERTEXT_WIDTH'd14315893;
publickey_row[4103] = `CIPHERTEXT_WIDTH'd5335067;
publickey_row[4104] = `CIPHERTEXT_WIDTH'd6651750;
publickey_row[4105] = `CIPHERTEXT_WIDTH'd929347;
publickey_row[4106] = `CIPHERTEXT_WIDTH'd12875625;
publickey_row[4107] = `CIPHERTEXT_WIDTH'd3985310;
publickey_row[4108] = `CIPHERTEXT_WIDTH'd12118107;
publickey_row[4109] = `CIPHERTEXT_WIDTH'd12950388;
publickey_row[4110] = `CIPHERTEXT_WIDTH'd358348;
publickey_row[4111] = `CIPHERTEXT_WIDTH'd16199464;
publickey_row[4112] = `CIPHERTEXT_WIDTH'd365246;
publickey_row[4113] = `CIPHERTEXT_WIDTH'd3186295;
publickey_row[4114] = `CIPHERTEXT_WIDTH'd11765324;
publickey_row[4115] = `CIPHERTEXT_WIDTH'd12028199;
publickey_row[4116] = `CIPHERTEXT_WIDTH'd15883183;
publickey_row[4117] = `CIPHERTEXT_WIDTH'd3291987;
publickey_row[4118] = `CIPHERTEXT_WIDTH'd3303834;
publickey_row[4119] = `CIPHERTEXT_WIDTH'd10477631;
publickey_row[4120] = `CIPHERTEXT_WIDTH'd6481055;
publickey_row[4121] = `CIPHERTEXT_WIDTH'd5925547;
publickey_row[4122] = `CIPHERTEXT_WIDTH'd7903289;
publickey_row[4123] = `CIPHERTEXT_WIDTH'd7383104;
publickey_row[4124] = `CIPHERTEXT_WIDTH'd9168427;
publickey_row[4125] = `CIPHERTEXT_WIDTH'd10166636;
publickey_row[4126] = `CIPHERTEXT_WIDTH'd8164985;
publickey_row[4127] = `CIPHERTEXT_WIDTH'd8173927;
publickey_row[4128] = `CIPHERTEXT_WIDTH'd14949261;
publickey_row[4129] = `CIPHERTEXT_WIDTH'd14244904;
publickey_row[4130] = `CIPHERTEXT_WIDTH'd7958185;
publickey_row[4131] = `CIPHERTEXT_WIDTH'd3743265;
publickey_row[4132] = `CIPHERTEXT_WIDTH'd1062255;
publickey_row[4133] = `CIPHERTEXT_WIDTH'd11151524;
publickey_row[4134] = `CIPHERTEXT_WIDTH'd1884627;
publickey_row[4135] = `CIPHERTEXT_WIDTH'd11049309;
publickey_row[4136] = `CIPHERTEXT_WIDTH'd6938770;
publickey_row[4137] = `CIPHERTEXT_WIDTH'd4602000;
publickey_row[4138] = `CIPHERTEXT_WIDTH'd16090530;
publickey_row[4139] = `CIPHERTEXT_WIDTH'd10248220;
publickey_row[4140] = `CIPHERTEXT_WIDTH'd8204853;
publickey_row[4141] = `CIPHERTEXT_WIDTH'd8493697;
publickey_row[4142] = `CIPHERTEXT_WIDTH'd14890711;
publickey_row[4143] = `CIPHERTEXT_WIDTH'd11185041;
publickey_row[4144] = `CIPHERTEXT_WIDTH'd10378763;
publickey_row[4145] = `CIPHERTEXT_WIDTH'd13931634;
publickey_row[4146] = `CIPHERTEXT_WIDTH'd4861632;
publickey_row[4147] = `CIPHERTEXT_WIDTH'd11867869;
publickey_row[4148] = `CIPHERTEXT_WIDTH'd10305413;
publickey_row[4149] = `CIPHERTEXT_WIDTH'd16059806;
publickey_row[4150] = `CIPHERTEXT_WIDTH'd5651964;
publickey_row[4151] = `CIPHERTEXT_WIDTH'd1671114;
publickey_row[4152] = `CIPHERTEXT_WIDTH'd3050157;
publickey_row[4153] = `CIPHERTEXT_WIDTH'd5517505;
publickey_row[4154] = `CIPHERTEXT_WIDTH'd15847415;
publickey_row[4155] = `CIPHERTEXT_WIDTH'd12988386;
publickey_row[4156] = `CIPHERTEXT_WIDTH'd8403667;
publickey_row[4157] = `CIPHERTEXT_WIDTH'd3871558;
publickey_row[4158] = `CIPHERTEXT_WIDTH'd8605692;
publickey_row[4159] = `CIPHERTEXT_WIDTH'd11560337;
publickey_row[4160] = `CIPHERTEXT_WIDTH'd8846779;
publickey_row[4161] = `CIPHERTEXT_WIDTH'd4582199;
publickey_row[4162] = `CIPHERTEXT_WIDTH'd7525241;
publickey_row[4163] = `CIPHERTEXT_WIDTH'd5036613;
publickey_row[4164] = `CIPHERTEXT_WIDTH'd8996687;
publickey_row[4165] = `CIPHERTEXT_WIDTH'd1782516;
publickey_row[4166] = `CIPHERTEXT_WIDTH'd10566042;
publickey_row[4167] = `CIPHERTEXT_WIDTH'd6643954;
publickey_row[4168] = `CIPHERTEXT_WIDTH'd10174995;
publickey_row[4169] = `CIPHERTEXT_WIDTH'd4868013;
publickey_row[4170] = `CIPHERTEXT_WIDTH'd9464892;
publickey_row[4171] = `CIPHERTEXT_WIDTH'd10827168;
publickey_row[4172] = `CIPHERTEXT_WIDTH'd1994063;
publickey_row[4173] = `CIPHERTEXT_WIDTH'd15610566;
publickey_row[4174] = `CIPHERTEXT_WIDTH'd7588002;
publickey_row[4175] = `CIPHERTEXT_WIDTH'd4847039;
publickey_row[4176] = `CIPHERTEXT_WIDTH'd3393862;
publickey_row[4177] = `CIPHERTEXT_WIDTH'd8587596;
publickey_row[4178] = `CIPHERTEXT_WIDTH'd14139597;
publickey_row[4179] = `CIPHERTEXT_WIDTH'd2241625;
publickey_row[4180] = `CIPHERTEXT_WIDTH'd2513794;
publickey_row[4181] = `CIPHERTEXT_WIDTH'd6062096;
publickey_row[4182] = `CIPHERTEXT_WIDTH'd238739;
publickey_row[4183] = `CIPHERTEXT_WIDTH'd14535934;
publickey_row[4184] = `CIPHERTEXT_WIDTH'd9339422;
publickey_row[4185] = `CIPHERTEXT_WIDTH'd4731502;
publickey_row[4186] = `CIPHERTEXT_WIDTH'd6938932;
publickey_row[4187] = `CIPHERTEXT_WIDTH'd1037996;
publickey_row[4188] = `CIPHERTEXT_WIDTH'd1263184;
publickey_row[4189] = `CIPHERTEXT_WIDTH'd7163763;
publickey_row[4190] = `CIPHERTEXT_WIDTH'd657330;
publickey_row[4191] = `CIPHERTEXT_WIDTH'd6411110;
publickey_row[4192] = `CIPHERTEXT_WIDTH'd14979499;
publickey_row[4193] = `CIPHERTEXT_WIDTH'd11506588;
publickey_row[4194] = `CIPHERTEXT_WIDTH'd144387;
publickey_row[4195] = `CIPHERTEXT_WIDTH'd6820017;
publickey_row[4196] = `CIPHERTEXT_WIDTH'd10423073;
publickey_row[4197] = `CIPHERTEXT_WIDTH'd8414408;
publickey_row[4198] = `CIPHERTEXT_WIDTH'd2566089;
publickey_row[4199] = `CIPHERTEXT_WIDTH'd8641868;
publickey_row[4200] = `CIPHERTEXT_WIDTH'd12474400;
publickey_row[4201] = `CIPHERTEXT_WIDTH'd1110132;
publickey_row[4202] = `CIPHERTEXT_WIDTH'd9071930;
publickey_row[4203] = `CIPHERTEXT_WIDTH'd5674177;
publickey_row[4204] = `CIPHERTEXT_WIDTH'd6532687;
publickey_row[4205] = `CIPHERTEXT_WIDTH'd4517829;
publickey_row[4206] = `CIPHERTEXT_WIDTH'd11511504;
publickey_row[4207] = `CIPHERTEXT_WIDTH'd5725102;
publickey_row[4208] = `CIPHERTEXT_WIDTH'd9405130;
publickey_row[4209] = `CIPHERTEXT_WIDTH'd4529403;
publickey_row[4210] = `CIPHERTEXT_WIDTH'd13266290;
publickey_row[4211] = `CIPHERTEXT_WIDTH'd9643876;
publickey_row[4212] = `CIPHERTEXT_WIDTH'd16082126;
publickey_row[4213] = `CIPHERTEXT_WIDTH'd7177145;
publickey_row[4214] = `CIPHERTEXT_WIDTH'd13075928;
publickey_row[4215] = `CIPHERTEXT_WIDTH'd12115786;
publickey_row[4216] = `CIPHERTEXT_WIDTH'd1433231;
publickey_row[4217] = `CIPHERTEXT_WIDTH'd4317721;
publickey_row[4218] = `CIPHERTEXT_WIDTH'd15459;
publickey_row[4219] = `CIPHERTEXT_WIDTH'd9455849;
publickey_row[4220] = `CIPHERTEXT_WIDTH'd16285049;
publickey_row[4221] = `CIPHERTEXT_WIDTH'd4740052;
publickey_row[4222] = `CIPHERTEXT_WIDTH'd761623;
publickey_row[4223] = `CIPHERTEXT_WIDTH'd99084;
publickey_row[4224] = `CIPHERTEXT_WIDTH'd3871681;
publickey_row[4225] = `CIPHERTEXT_WIDTH'd6908275;
publickey_row[4226] = `CIPHERTEXT_WIDTH'd4240509;
publickey_row[4227] = `CIPHERTEXT_WIDTH'd11678444;
publickey_row[4228] = `CIPHERTEXT_WIDTH'd3840920;
publickey_row[4229] = `CIPHERTEXT_WIDTH'd2404588;
publickey_row[4230] = `CIPHERTEXT_WIDTH'd11435020;
publickey_row[4231] = `CIPHERTEXT_WIDTH'd13981276;
publickey_row[4232] = `CIPHERTEXT_WIDTH'd7869558;
publickey_row[4233] = `CIPHERTEXT_WIDTH'd10963310;
publickey_row[4234] = `CIPHERTEXT_WIDTH'd15709686;
publickey_row[4235] = `CIPHERTEXT_WIDTH'd665714;
publickey_row[4236] = `CIPHERTEXT_WIDTH'd8512798;
publickey_row[4237] = `CIPHERTEXT_WIDTH'd10486757;
publickey_row[4238] = `CIPHERTEXT_WIDTH'd3524383;
publickey_row[4239] = `CIPHERTEXT_WIDTH'd11847405;
publickey_row[4240] = `CIPHERTEXT_WIDTH'd4329330;
publickey_row[4241] = `CIPHERTEXT_WIDTH'd6515478;
publickey_row[4242] = `CIPHERTEXT_WIDTH'd16279340;
publickey_row[4243] = `CIPHERTEXT_WIDTH'd13139381;
publickey_row[4244] = `CIPHERTEXT_WIDTH'd11239729;
publickey_row[4245] = `CIPHERTEXT_WIDTH'd4643660;
publickey_row[4246] = `CIPHERTEXT_WIDTH'd14081476;
publickey_row[4247] = `CIPHERTEXT_WIDTH'd7831552;
publickey_row[4248] = `CIPHERTEXT_WIDTH'd101867;
publickey_row[4249] = `CIPHERTEXT_WIDTH'd16277118;
publickey_row[4250] = `CIPHERTEXT_WIDTH'd12951267;
publickey_row[4251] = `CIPHERTEXT_WIDTH'd13375038;
publickey_row[4252] = `CIPHERTEXT_WIDTH'd211802;
publickey_row[4253] = `CIPHERTEXT_WIDTH'd7455007;
publickey_row[4254] = `CIPHERTEXT_WIDTH'd3845179;
publickey_row[4255] = `CIPHERTEXT_WIDTH'd1130915;
publickey_row[4256] = `CIPHERTEXT_WIDTH'd5871215;
publickey_row[4257] = `CIPHERTEXT_WIDTH'd11591356;
publickey_row[4258] = `CIPHERTEXT_WIDTH'd15261347;
publickey_row[4259] = `CIPHERTEXT_WIDTH'd13362207;
publickey_row[4260] = `CIPHERTEXT_WIDTH'd12835499;
publickey_row[4261] = `CIPHERTEXT_WIDTH'd7774887;
publickey_row[4262] = `CIPHERTEXT_WIDTH'd14179468;
publickey_row[4263] = `CIPHERTEXT_WIDTH'd7564344;
publickey_row[4264] = `CIPHERTEXT_WIDTH'd899985;
publickey_row[4265] = `CIPHERTEXT_WIDTH'd4840710;
publickey_row[4266] = `CIPHERTEXT_WIDTH'd10665287;
publickey_row[4267] = `CIPHERTEXT_WIDTH'd7439035;
publickey_row[4268] = `CIPHERTEXT_WIDTH'd9303691;
publickey_row[4269] = `CIPHERTEXT_WIDTH'd8550792;
publickey_row[4270] = `CIPHERTEXT_WIDTH'd14835371;
publickey_row[4271] = `CIPHERTEXT_WIDTH'd8332351;
publickey_row[4272] = `CIPHERTEXT_WIDTH'd7084499;
publickey_row[4273] = `CIPHERTEXT_WIDTH'd13682930;
publickey_row[4274] = `CIPHERTEXT_WIDTH'd4570837;
publickey_row[4275] = `CIPHERTEXT_WIDTH'd10990796;
publickey_row[4276] = `CIPHERTEXT_WIDTH'd12318225;
publickey_row[4277] = `CIPHERTEXT_WIDTH'd2832278;
publickey_row[4278] = `CIPHERTEXT_WIDTH'd15592688;
publickey_row[4279] = `CIPHERTEXT_WIDTH'd12760544;
publickey_row[4280] = `CIPHERTEXT_WIDTH'd15337130;
publickey_row[4281] = `CIPHERTEXT_WIDTH'd11656267;
publickey_row[4282] = `CIPHERTEXT_WIDTH'd14105084;
publickey_row[4283] = `CIPHERTEXT_WIDTH'd10783339;
publickey_row[4284] = `CIPHERTEXT_WIDTH'd9862207;
publickey_row[4285] = `CIPHERTEXT_WIDTH'd14735448;
publickey_row[4286] = `CIPHERTEXT_WIDTH'd3277770;
publickey_row[4287] = `CIPHERTEXT_WIDTH'd11556096;
publickey_row[4288] = `CIPHERTEXT_WIDTH'd10729532;
publickey_row[4289] = `CIPHERTEXT_WIDTH'd4897054;
publickey_row[4290] = `CIPHERTEXT_WIDTH'd8942525;
publickey_row[4291] = `CIPHERTEXT_WIDTH'd14966258;
publickey_row[4292] = `CIPHERTEXT_WIDTH'd3378428;
publickey_row[4293] = `CIPHERTEXT_WIDTH'd2705316;
publickey_row[4294] = `CIPHERTEXT_WIDTH'd13263016;
publickey_row[4295] = `CIPHERTEXT_WIDTH'd7514898;
publickey_row[4296] = `CIPHERTEXT_WIDTH'd10347818;
publickey_row[4297] = `CIPHERTEXT_WIDTH'd10310750;
publickey_row[4298] = `CIPHERTEXT_WIDTH'd9343639;
publickey_row[4299] = `CIPHERTEXT_WIDTH'd16408848;
publickey_row[4300] = `CIPHERTEXT_WIDTH'd15603733;
publickey_row[4301] = `CIPHERTEXT_WIDTH'd11620309;
publickey_row[4302] = `CIPHERTEXT_WIDTH'd14771202;
publickey_row[4303] = `CIPHERTEXT_WIDTH'd15610421;
publickey_row[4304] = `CIPHERTEXT_WIDTH'd4108616;
publickey_row[4305] = `CIPHERTEXT_WIDTH'd5531522;
publickey_row[4306] = `CIPHERTEXT_WIDTH'd9494303;
publickey_row[4307] = `CIPHERTEXT_WIDTH'd5153723;
publickey_row[4308] = `CIPHERTEXT_WIDTH'd7689510;
publickey_row[4309] = `CIPHERTEXT_WIDTH'd3953064;
publickey_row[4310] = `CIPHERTEXT_WIDTH'd15209018;
publickey_row[4311] = `CIPHERTEXT_WIDTH'd13448751;
publickey_row[4312] = `CIPHERTEXT_WIDTH'd12844656;
publickey_row[4313] = `CIPHERTEXT_WIDTH'd14168662;
publickey_row[4314] = `CIPHERTEXT_WIDTH'd6853582;
publickey_row[4315] = `CIPHERTEXT_WIDTH'd4047451;
publickey_row[4316] = `CIPHERTEXT_WIDTH'd10649605;
publickey_row[4317] = `CIPHERTEXT_WIDTH'd12020600;
publickey_row[4318] = `CIPHERTEXT_WIDTH'd5468877;
publickey_row[4319] = `CIPHERTEXT_WIDTH'd14380141;
publickey_row[4320] = `CIPHERTEXT_WIDTH'd13533935;
publickey_row[4321] = `CIPHERTEXT_WIDTH'd13528002;
publickey_row[4322] = `CIPHERTEXT_WIDTH'd13378991;
publickey_row[4323] = `CIPHERTEXT_WIDTH'd13796743;
publickey_row[4324] = `CIPHERTEXT_WIDTH'd15225303;
publickey_row[4325] = `CIPHERTEXT_WIDTH'd15502855;
publickey_row[4326] = `CIPHERTEXT_WIDTH'd8104945;
publickey_row[4327] = `CIPHERTEXT_WIDTH'd13508910;
publickey_row[4328] = `CIPHERTEXT_WIDTH'd11653031;
publickey_row[4329] = `CIPHERTEXT_WIDTH'd13509806;
publickey_row[4330] = `CIPHERTEXT_WIDTH'd8828802;
publickey_row[4331] = `CIPHERTEXT_WIDTH'd311492;
publickey_row[4332] = `CIPHERTEXT_WIDTH'd3023823;
publickey_row[4333] = `CIPHERTEXT_WIDTH'd3082162;
publickey_row[4334] = `CIPHERTEXT_WIDTH'd13439648;
publickey_row[4335] = `CIPHERTEXT_WIDTH'd1975217;
publickey_row[4336] = `CIPHERTEXT_WIDTH'd7541465;
publickey_row[4337] = `CIPHERTEXT_WIDTH'd1857300;
publickey_row[4338] = `CIPHERTEXT_WIDTH'd844245;
publickey_row[4339] = `CIPHERTEXT_WIDTH'd5370912;
publickey_row[4340] = `CIPHERTEXT_WIDTH'd8604914;
publickey_row[4341] = `CIPHERTEXT_WIDTH'd3034555;
publickey_row[4342] = `CIPHERTEXT_WIDTH'd6969424;
publickey_row[4343] = `CIPHERTEXT_WIDTH'd14441778;
publickey_row[4344] = `CIPHERTEXT_WIDTH'd7101990;
publickey_row[4345] = `CIPHERTEXT_WIDTH'd5577251;
publickey_row[4346] = `CIPHERTEXT_WIDTH'd8027536;
publickey_row[4347] = `CIPHERTEXT_WIDTH'd11936962;
publickey_row[4348] = `CIPHERTEXT_WIDTH'd5657259;
publickey_row[4349] = `CIPHERTEXT_WIDTH'd7629270;
publickey_row[4350] = `CIPHERTEXT_WIDTH'd11351088;
publickey_row[4351] = `CIPHERTEXT_WIDTH'd192063;
publickey_row[4352] = `CIPHERTEXT_WIDTH'd15422556;
publickey_row[4353] = `CIPHERTEXT_WIDTH'd7785010;
publickey_row[4354] = `CIPHERTEXT_WIDTH'd8664468;
publickey_row[4355] = `CIPHERTEXT_WIDTH'd8818069;
publickey_row[4356] = `CIPHERTEXT_WIDTH'd4305715;
publickey_row[4357] = `CIPHERTEXT_WIDTH'd1642773;
publickey_row[4358] = `CIPHERTEXT_WIDTH'd6299737;
publickey_row[4359] = `CIPHERTEXT_WIDTH'd1404508;
publickey_row[4360] = `CIPHERTEXT_WIDTH'd14264149;
publickey_row[4361] = `CIPHERTEXT_WIDTH'd251539;
publickey_row[4362] = `CIPHERTEXT_WIDTH'd11186588;
publickey_row[4363] = `CIPHERTEXT_WIDTH'd13981575;
publickey_row[4364] = `CIPHERTEXT_WIDTH'd4198033;
publickey_row[4365] = `CIPHERTEXT_WIDTH'd6535266;
publickey_row[4366] = `CIPHERTEXT_WIDTH'd521976;
publickey_row[4367] = `CIPHERTEXT_WIDTH'd14527680;
publickey_row[4368] = `CIPHERTEXT_WIDTH'd12402563;
publickey_row[4369] = `CIPHERTEXT_WIDTH'd16233590;
publickey_row[4370] = `CIPHERTEXT_WIDTH'd950432;
publickey_row[4371] = `CIPHERTEXT_WIDTH'd13667977;
publickey_row[4372] = `CIPHERTEXT_WIDTH'd937152;
publickey_row[4373] = `CIPHERTEXT_WIDTH'd5632680;
publickey_row[4374] = `CIPHERTEXT_WIDTH'd12730964;
publickey_row[4375] = `CIPHERTEXT_WIDTH'd552331;
publickey_row[4376] = `CIPHERTEXT_WIDTH'd9804181;
publickey_row[4377] = `CIPHERTEXT_WIDTH'd1256005;
publickey_row[4378] = `CIPHERTEXT_WIDTH'd5691097;
publickey_row[4379] = `CIPHERTEXT_WIDTH'd13366831;
publickey_row[4380] = `CIPHERTEXT_WIDTH'd16321461;
publickey_row[4381] = `CIPHERTEXT_WIDTH'd7866351;
publickey_row[4382] = `CIPHERTEXT_WIDTH'd1902482;
publickey_row[4383] = `CIPHERTEXT_WIDTH'd10868646;
publickey_row[4384] = `CIPHERTEXT_WIDTH'd7134676;
publickey_row[4385] = `CIPHERTEXT_WIDTH'd2145417;
publickey_row[4386] = `CIPHERTEXT_WIDTH'd3746294;
publickey_row[4387] = `CIPHERTEXT_WIDTH'd936503;
publickey_row[4388] = `CIPHERTEXT_WIDTH'd2913469;
publickey_row[4389] = `CIPHERTEXT_WIDTH'd3082768;
publickey_row[4390] = `CIPHERTEXT_WIDTH'd9105014;
publickey_row[4391] = `CIPHERTEXT_WIDTH'd701809;
publickey_row[4392] = `CIPHERTEXT_WIDTH'd16417720;
publickey_row[4393] = `CIPHERTEXT_WIDTH'd14884301;
publickey_row[4394] = `CIPHERTEXT_WIDTH'd8844764;
publickey_row[4395] = `CIPHERTEXT_WIDTH'd12191239;
publickey_row[4396] = `CIPHERTEXT_WIDTH'd6634631;
publickey_row[4397] = `CIPHERTEXT_WIDTH'd7741526;
publickey_row[4398] = `CIPHERTEXT_WIDTH'd16315970;
publickey_row[4399] = `CIPHERTEXT_WIDTH'd4915458;
publickey_row[4400] = `CIPHERTEXT_WIDTH'd6367199;
publickey_row[4401] = `CIPHERTEXT_WIDTH'd8419127;
publickey_row[4402] = `CIPHERTEXT_WIDTH'd5812795;
publickey_row[4403] = `CIPHERTEXT_WIDTH'd3095041;
publickey_row[4404] = `CIPHERTEXT_WIDTH'd846236;
publickey_row[4405] = `CIPHERTEXT_WIDTH'd6301898;
publickey_row[4406] = `CIPHERTEXT_WIDTH'd2753245;
publickey_row[4407] = `CIPHERTEXT_WIDTH'd16655585;
publickey_row[4408] = `CIPHERTEXT_WIDTH'd11378946;
publickey_row[4409] = `CIPHERTEXT_WIDTH'd5647845;
publickey_row[4410] = `CIPHERTEXT_WIDTH'd4013000;
publickey_row[4411] = `CIPHERTEXT_WIDTH'd11439074;
publickey_row[4412] = `CIPHERTEXT_WIDTH'd3938423;
publickey_row[4413] = `CIPHERTEXT_WIDTH'd12511682;
publickey_row[4414] = `CIPHERTEXT_WIDTH'd4982835;
publickey_row[4415] = `CIPHERTEXT_WIDTH'd11230936;
publickey_row[4416] = `CIPHERTEXT_WIDTH'd10751135;
publickey_row[4417] = `CIPHERTEXT_WIDTH'd4892643;
publickey_row[4418] = `CIPHERTEXT_WIDTH'd11868097;
publickey_row[4419] = `CIPHERTEXT_WIDTH'd992375;
publickey_row[4420] = `CIPHERTEXT_WIDTH'd8496486;
publickey_row[4421] = `CIPHERTEXT_WIDTH'd12512644;
publickey_row[4422] = `CIPHERTEXT_WIDTH'd4400961;
publickey_row[4423] = `CIPHERTEXT_WIDTH'd4820327;
publickey_row[4424] = `CIPHERTEXT_WIDTH'd6837335;
publickey_row[4425] = `CIPHERTEXT_WIDTH'd4055410;
publickey_row[4426] = `CIPHERTEXT_WIDTH'd8005765;
publickey_row[4427] = `CIPHERTEXT_WIDTH'd15188376;
publickey_row[4428] = `CIPHERTEXT_WIDTH'd15837546;
publickey_row[4429] = `CIPHERTEXT_WIDTH'd4347475;
publickey_row[4430] = `CIPHERTEXT_WIDTH'd3404389;
publickey_row[4431] = `CIPHERTEXT_WIDTH'd9088045;
publickey_row[4432] = `CIPHERTEXT_WIDTH'd11960099;
publickey_row[4433] = `CIPHERTEXT_WIDTH'd2920837;
publickey_row[4434] = `CIPHERTEXT_WIDTH'd1810033;
publickey_row[4435] = `CIPHERTEXT_WIDTH'd4135449;
publickey_row[4436] = `CIPHERTEXT_WIDTH'd1880154;
publickey_row[4437] = `CIPHERTEXT_WIDTH'd14755671;
publickey_row[4438] = `CIPHERTEXT_WIDTH'd9865515;
publickey_row[4439] = `CIPHERTEXT_WIDTH'd794390;
publickey_row[4440] = `CIPHERTEXT_WIDTH'd16067771;
publickey_row[4441] = `CIPHERTEXT_WIDTH'd1603135;
publickey_row[4442] = `CIPHERTEXT_WIDTH'd13802451;
publickey_row[4443] = `CIPHERTEXT_WIDTH'd15374393;
publickey_row[4444] = `CIPHERTEXT_WIDTH'd10869654;
publickey_row[4445] = `CIPHERTEXT_WIDTH'd14725671;
publickey_row[4446] = `CIPHERTEXT_WIDTH'd12062456;
publickey_row[4447] = `CIPHERTEXT_WIDTH'd14224879;
publickey_row[4448] = `CIPHERTEXT_WIDTH'd11957200;
publickey_row[4449] = `CIPHERTEXT_WIDTH'd10429663;
publickey_row[4450] = `CIPHERTEXT_WIDTH'd11434436;
publickey_row[4451] = `CIPHERTEXT_WIDTH'd3453882;
publickey_row[4452] = `CIPHERTEXT_WIDTH'd11608609;
publickey_row[4453] = `CIPHERTEXT_WIDTH'd2111930;
publickey_row[4454] = `CIPHERTEXT_WIDTH'd2726892;
publickey_row[4455] = `CIPHERTEXT_WIDTH'd3214132;
publickey_row[4456] = `CIPHERTEXT_WIDTH'd16262976;
publickey_row[4457] = `CIPHERTEXT_WIDTH'd1441691;
publickey_row[4458] = `CIPHERTEXT_WIDTH'd12696011;
publickey_row[4459] = `CIPHERTEXT_WIDTH'd10819944;
publickey_row[4460] = `CIPHERTEXT_WIDTH'd14096637;
publickey_row[4461] = `CIPHERTEXT_WIDTH'd2400350;
publickey_row[4462] = `CIPHERTEXT_WIDTH'd4484482;
publickey_row[4463] = `CIPHERTEXT_WIDTH'd3485253;
publickey_row[4464] = `CIPHERTEXT_WIDTH'd4151494;
publickey_row[4465] = `CIPHERTEXT_WIDTH'd15049165;
publickey_row[4466] = `CIPHERTEXT_WIDTH'd109756;
publickey_row[4467] = `CIPHERTEXT_WIDTH'd2680763;
publickey_row[4468] = `CIPHERTEXT_WIDTH'd14328476;
publickey_row[4469] = `CIPHERTEXT_WIDTH'd16520568;
publickey_row[4470] = `CIPHERTEXT_WIDTH'd585084;
publickey_row[4471] = `CIPHERTEXT_WIDTH'd10190984;
publickey_row[4472] = `CIPHERTEXT_WIDTH'd9742760;
publickey_row[4473] = `CIPHERTEXT_WIDTH'd4460790;
publickey_row[4474] = `CIPHERTEXT_WIDTH'd6979100;
publickey_row[4475] = `CIPHERTEXT_WIDTH'd7171660;
publickey_row[4476] = `CIPHERTEXT_WIDTH'd5539275;
publickey_row[4477] = `CIPHERTEXT_WIDTH'd5888936;
publickey_row[4478] = `CIPHERTEXT_WIDTH'd15614183;
publickey_row[4479] = `CIPHERTEXT_WIDTH'd808693;
publickey_row[4480] = `CIPHERTEXT_WIDTH'd5336987;
publickey_row[4481] = `CIPHERTEXT_WIDTH'd11105369;
publickey_row[4482] = `CIPHERTEXT_WIDTH'd13556057;
publickey_row[4483] = `CIPHERTEXT_WIDTH'd9475767;
publickey_row[4484] = `CIPHERTEXT_WIDTH'd14884165;
publickey_row[4485] = `CIPHERTEXT_WIDTH'd15730050;
publickey_row[4486] = `CIPHERTEXT_WIDTH'd3859083;
publickey_row[4487] = `CIPHERTEXT_WIDTH'd12692456;
publickey_row[4488] = `CIPHERTEXT_WIDTH'd2894177;
publickey_row[4489] = `CIPHERTEXT_WIDTH'd7735795;
publickey_row[4490] = `CIPHERTEXT_WIDTH'd10690530;
publickey_row[4491] = `CIPHERTEXT_WIDTH'd1179533;
publickey_row[4492] = `CIPHERTEXT_WIDTH'd5492835;
publickey_row[4493] = `CIPHERTEXT_WIDTH'd1559665;
publickey_row[4494] = `CIPHERTEXT_WIDTH'd10270027;
publickey_row[4495] = `CIPHERTEXT_WIDTH'd13594772;
publickey_row[4496] = `CIPHERTEXT_WIDTH'd5051911;
publickey_row[4497] = `CIPHERTEXT_WIDTH'd6586667;
publickey_row[4498] = `CIPHERTEXT_WIDTH'd10707269;
publickey_row[4499] = `CIPHERTEXT_WIDTH'd9049750;
publickey_row[4500] = `CIPHERTEXT_WIDTH'd7228541;
publickey_row[4501] = `CIPHERTEXT_WIDTH'd6401593;
publickey_row[4502] = `CIPHERTEXT_WIDTH'd15298207;
publickey_row[4503] = `CIPHERTEXT_WIDTH'd275848;
publickey_row[4504] = `CIPHERTEXT_WIDTH'd14787705;
publickey_row[4505] = `CIPHERTEXT_WIDTH'd1403593;
publickey_row[4506] = `CIPHERTEXT_WIDTH'd1897689;
publickey_row[4507] = `CIPHERTEXT_WIDTH'd15869971;
publickey_row[4508] = `CIPHERTEXT_WIDTH'd4081783;
publickey_row[4509] = `CIPHERTEXT_WIDTH'd11904548;
publickey_row[4510] = `CIPHERTEXT_WIDTH'd3889219;
publickey_row[4511] = `CIPHERTEXT_WIDTH'd9793250;
publickey_row[4512] = `CIPHERTEXT_WIDTH'd2296703;
publickey_row[4513] = `CIPHERTEXT_WIDTH'd3627892;
publickey_row[4514] = `CIPHERTEXT_WIDTH'd14426482;
publickey_row[4515] = `CIPHERTEXT_WIDTH'd9068660;
publickey_row[4516] = `CIPHERTEXT_WIDTH'd4002987;
publickey_row[4517] = `CIPHERTEXT_WIDTH'd9650746;
publickey_row[4518] = `CIPHERTEXT_WIDTH'd1985845;
publickey_row[4519] = `CIPHERTEXT_WIDTH'd6644788;
publickey_row[4520] = `CIPHERTEXT_WIDTH'd8792259;
publickey_row[4521] = `CIPHERTEXT_WIDTH'd14186327;
publickey_row[4522] = `CIPHERTEXT_WIDTH'd2596334;
publickey_row[4523] = `CIPHERTEXT_WIDTH'd12206443;
publickey_row[4524] = `CIPHERTEXT_WIDTH'd3969396;
publickey_row[4525] = `CIPHERTEXT_WIDTH'd11081990;
publickey_row[4526] = `CIPHERTEXT_WIDTH'd15518103;
publickey_row[4527] = `CIPHERTEXT_WIDTH'd3267489;
publickey_row[4528] = `CIPHERTEXT_WIDTH'd401617;
publickey_row[4529] = `CIPHERTEXT_WIDTH'd13020827;
publickey_row[4530] = `CIPHERTEXT_WIDTH'd11912639;
publickey_row[4531] = `CIPHERTEXT_WIDTH'd5513160;
publickey_row[4532] = `CIPHERTEXT_WIDTH'd15455766;
publickey_row[4533] = `CIPHERTEXT_WIDTH'd10160921;
publickey_row[4534] = `CIPHERTEXT_WIDTH'd15203417;
publickey_row[4535] = `CIPHERTEXT_WIDTH'd12215113;
publickey_row[4536] = `CIPHERTEXT_WIDTH'd5247960;
publickey_row[4537] = `CIPHERTEXT_WIDTH'd2141612;
publickey_row[4538] = `CIPHERTEXT_WIDTH'd15430142;
publickey_row[4539] = `CIPHERTEXT_WIDTH'd5276795;
publickey_row[4540] = `CIPHERTEXT_WIDTH'd9882987;
publickey_row[4541] = `CIPHERTEXT_WIDTH'd5253131;
publickey_row[4542] = `CIPHERTEXT_WIDTH'd5335622;
publickey_row[4543] = `CIPHERTEXT_WIDTH'd1937694;
publickey_row[4544] = `CIPHERTEXT_WIDTH'd14568596;
publickey_row[4545] = `CIPHERTEXT_WIDTH'd4982738;
publickey_row[4546] = `CIPHERTEXT_WIDTH'd13631112;
publickey_row[4547] = `CIPHERTEXT_WIDTH'd1675977;
publickey_row[4548] = `CIPHERTEXT_WIDTH'd8461566;
publickey_row[4549] = `CIPHERTEXT_WIDTH'd13808011;
publickey_row[4550] = `CIPHERTEXT_WIDTH'd6640139;
publickey_row[4551] = `CIPHERTEXT_WIDTH'd3130544;
publickey_row[4552] = `CIPHERTEXT_WIDTH'd6742696;
publickey_row[4553] = `CIPHERTEXT_WIDTH'd8154751;
publickey_row[4554] = `CIPHERTEXT_WIDTH'd10267583;
publickey_row[4555] = `CIPHERTEXT_WIDTH'd11728099;
publickey_row[4556] = `CIPHERTEXT_WIDTH'd4328461;
publickey_row[4557] = `CIPHERTEXT_WIDTH'd10760468;
publickey_row[4558] = `CIPHERTEXT_WIDTH'd4513774;
publickey_row[4559] = `CIPHERTEXT_WIDTH'd221335;
publickey_row[4560] = `CIPHERTEXT_WIDTH'd4130731;
publickey_row[4561] = `CIPHERTEXT_WIDTH'd11710792;
publickey_row[4562] = `CIPHERTEXT_WIDTH'd16267998;
publickey_row[4563] = `CIPHERTEXT_WIDTH'd4358377;
publickey_row[4564] = `CIPHERTEXT_WIDTH'd2279526;
publickey_row[4565] = `CIPHERTEXT_WIDTH'd7959307;
publickey_row[4566] = `CIPHERTEXT_WIDTH'd5212534;
publickey_row[4567] = `CIPHERTEXT_WIDTH'd5285752;
publickey_row[4568] = `CIPHERTEXT_WIDTH'd10813595;
publickey_row[4569] = `CIPHERTEXT_WIDTH'd1793574;
publickey_row[4570] = `CIPHERTEXT_WIDTH'd6695000;
publickey_row[4571] = `CIPHERTEXT_WIDTH'd2398206;
publickey_row[4572] = `CIPHERTEXT_WIDTH'd8186777;
publickey_row[4573] = `CIPHERTEXT_WIDTH'd13497973;
publickey_row[4574] = `CIPHERTEXT_WIDTH'd1707298;
publickey_row[4575] = `CIPHERTEXT_WIDTH'd1596050;
publickey_row[4576] = `CIPHERTEXT_WIDTH'd10582049;
publickey_row[4577] = `CIPHERTEXT_WIDTH'd12431514;
publickey_row[4578] = `CIPHERTEXT_WIDTH'd6112378;
publickey_row[4579] = `CIPHERTEXT_WIDTH'd1769005;
publickey_row[4580] = `CIPHERTEXT_WIDTH'd13868471;
publickey_row[4581] = `CIPHERTEXT_WIDTH'd14806099;
publickey_row[4582] = `CIPHERTEXT_WIDTH'd14360137;
publickey_row[4583] = `CIPHERTEXT_WIDTH'd1194705;
publickey_row[4584] = `CIPHERTEXT_WIDTH'd2316339;
publickey_row[4585] = `CIPHERTEXT_WIDTH'd9766688;
publickey_row[4586] = `CIPHERTEXT_WIDTH'd4135492;
publickey_row[4587] = `CIPHERTEXT_WIDTH'd6601518;
publickey_row[4588] = `CIPHERTEXT_WIDTH'd4278661;
publickey_row[4589] = `CIPHERTEXT_WIDTH'd3379515;
publickey_row[4590] = `CIPHERTEXT_WIDTH'd5676735;
publickey_row[4591] = `CIPHERTEXT_WIDTH'd7905365;
publickey_row[4592] = `CIPHERTEXT_WIDTH'd1420184;
publickey_row[4593] = `CIPHERTEXT_WIDTH'd11713060;
publickey_row[4594] = `CIPHERTEXT_WIDTH'd4372232;
publickey_row[4595] = `CIPHERTEXT_WIDTH'd4368774;
publickey_row[4596] = `CIPHERTEXT_WIDTH'd6158299;
publickey_row[4597] = `CIPHERTEXT_WIDTH'd12300799;
publickey_row[4598] = `CIPHERTEXT_WIDTH'd11510088;
publickey_row[4599] = `CIPHERTEXT_WIDTH'd1360761;
publickey_row[4600] = `CIPHERTEXT_WIDTH'd16334831;
publickey_row[4601] = `CIPHERTEXT_WIDTH'd1257939;
publickey_row[4602] = `CIPHERTEXT_WIDTH'd7362517;
publickey_row[4603] = `CIPHERTEXT_WIDTH'd7736469;
publickey_row[4604] = `CIPHERTEXT_WIDTH'd676701;
publickey_row[4605] = `CIPHERTEXT_WIDTH'd2007677;
publickey_row[4606] = `CIPHERTEXT_WIDTH'd13673178;
publickey_row[4607] = `CIPHERTEXT_WIDTH'd16420134;
publickey_row[4608] = `CIPHERTEXT_WIDTH'd2012749;
publickey_row[4609] = `CIPHERTEXT_WIDTH'd13403663;
publickey_row[4610] = `CIPHERTEXT_WIDTH'd15962115;
publickey_row[4611] = `CIPHERTEXT_WIDTH'd5116354;
publickey_row[4612] = `CIPHERTEXT_WIDTH'd1864436;
publickey_row[4613] = `CIPHERTEXT_WIDTH'd9563512;
publickey_row[4614] = `CIPHERTEXT_WIDTH'd12388719;
publickey_row[4615] = `CIPHERTEXT_WIDTH'd12787444;
publickey_row[4616] = `CIPHERTEXT_WIDTH'd4191275;
publickey_row[4617] = `CIPHERTEXT_WIDTH'd6194830;
publickey_row[4618] = `CIPHERTEXT_WIDTH'd13261362;
publickey_row[4619] = `CIPHERTEXT_WIDTH'd1603608;
publickey_row[4620] = `CIPHERTEXT_WIDTH'd14335043;
publickey_row[4621] = `CIPHERTEXT_WIDTH'd5693410;
publickey_row[4622] = `CIPHERTEXT_WIDTH'd3285660;
publickey_row[4623] = `CIPHERTEXT_WIDTH'd12229231;
publickey_row[4624] = `CIPHERTEXT_WIDTH'd6916491;
publickey_row[4625] = `CIPHERTEXT_WIDTH'd2006307;
publickey_row[4626] = `CIPHERTEXT_WIDTH'd9231195;
publickey_row[4627] = `CIPHERTEXT_WIDTH'd14396467;
publickey_row[4628] = `CIPHERTEXT_WIDTH'd10056552;
publickey_row[4629] = `CIPHERTEXT_WIDTH'd12183203;
publickey_row[4630] = `CIPHERTEXT_WIDTH'd9746662;
publickey_row[4631] = `CIPHERTEXT_WIDTH'd15104777;
publickey_row[4632] = `CIPHERTEXT_WIDTH'd15569255;
publickey_row[4633] = `CIPHERTEXT_WIDTH'd8014234;
publickey_row[4634] = `CIPHERTEXT_WIDTH'd12752622;
publickey_row[4635] = `CIPHERTEXT_WIDTH'd2321381;
publickey_row[4636] = `CIPHERTEXT_WIDTH'd12263266;
publickey_row[4637] = `CIPHERTEXT_WIDTH'd4565976;
publickey_row[4638] = `CIPHERTEXT_WIDTH'd306951;
publickey_row[4639] = `CIPHERTEXT_WIDTH'd8598812;
publickey_row[4640] = `CIPHERTEXT_WIDTH'd12678616;
publickey_row[4641] = `CIPHERTEXT_WIDTH'd7526771;
publickey_row[4642] = `CIPHERTEXT_WIDTH'd1145824;
publickey_row[4643] = `CIPHERTEXT_WIDTH'd12982985;
publickey_row[4644] = `CIPHERTEXT_WIDTH'd4806101;
publickey_row[4645] = `CIPHERTEXT_WIDTH'd14915414;
publickey_row[4646] = `CIPHERTEXT_WIDTH'd6598979;
publickey_row[4647] = `CIPHERTEXT_WIDTH'd10919861;
publickey_row[4648] = `CIPHERTEXT_WIDTH'd9481452;
publickey_row[4649] = `CIPHERTEXT_WIDTH'd12722012;
publickey_row[4650] = `CIPHERTEXT_WIDTH'd13991585;
publickey_row[4651] = `CIPHERTEXT_WIDTH'd9123615;
publickey_row[4652] = `CIPHERTEXT_WIDTH'd5553325;
publickey_row[4653] = `CIPHERTEXT_WIDTH'd6763272;
publickey_row[4654] = `CIPHERTEXT_WIDTH'd9685896;
publickey_row[4655] = `CIPHERTEXT_WIDTH'd721094;
publickey_row[4656] = `CIPHERTEXT_WIDTH'd6581771;
publickey_row[4657] = `CIPHERTEXT_WIDTH'd13653307;
publickey_row[4658] = `CIPHERTEXT_WIDTH'd12947851;
publickey_row[4659] = `CIPHERTEXT_WIDTH'd9702498;
publickey_row[4660] = `CIPHERTEXT_WIDTH'd12728168;
publickey_row[4661] = `CIPHERTEXT_WIDTH'd4378793;
publickey_row[4662] = `CIPHERTEXT_WIDTH'd8552761;
publickey_row[4663] = `CIPHERTEXT_WIDTH'd233711;
publickey_row[4664] = `CIPHERTEXT_WIDTH'd7919456;
publickey_row[4665] = `CIPHERTEXT_WIDTH'd9644666;
publickey_row[4666] = `CIPHERTEXT_WIDTH'd7848813;
publickey_row[4667] = `CIPHERTEXT_WIDTH'd3825038;
publickey_row[4668] = `CIPHERTEXT_WIDTH'd1655747;
publickey_row[4669] = `CIPHERTEXT_WIDTH'd11916566;
publickey_row[4670] = `CIPHERTEXT_WIDTH'd2704807;
publickey_row[4671] = `CIPHERTEXT_WIDTH'd10445738;
publickey_row[4672] = `CIPHERTEXT_WIDTH'd5809117;
publickey_row[4673] = `CIPHERTEXT_WIDTH'd3565179;
publickey_row[4674] = `CIPHERTEXT_WIDTH'd15661935;
publickey_row[4675] = `CIPHERTEXT_WIDTH'd16527025;
publickey_row[4676] = `CIPHERTEXT_WIDTH'd16097990;
publickey_row[4677] = `CIPHERTEXT_WIDTH'd16760510;
publickey_row[4678] = `CIPHERTEXT_WIDTH'd6038619;
publickey_row[4679] = `CIPHERTEXT_WIDTH'd5807505;
publickey_row[4680] = `CIPHERTEXT_WIDTH'd3606941;
publickey_row[4681] = `CIPHERTEXT_WIDTH'd10626510;
publickey_row[4682] = `CIPHERTEXT_WIDTH'd8655431;
publickey_row[4683] = `CIPHERTEXT_WIDTH'd7203345;
publickey_row[4684] = `CIPHERTEXT_WIDTH'd1225064;
publickey_row[4685] = `CIPHERTEXT_WIDTH'd14851079;
publickey_row[4686] = `CIPHERTEXT_WIDTH'd3494612;
publickey_row[4687] = `CIPHERTEXT_WIDTH'd6117576;
publickey_row[4688] = `CIPHERTEXT_WIDTH'd2671078;
publickey_row[4689] = `CIPHERTEXT_WIDTH'd15346372;
publickey_row[4690] = `CIPHERTEXT_WIDTH'd9849025;
publickey_row[4691] = `CIPHERTEXT_WIDTH'd2753698;
publickey_row[4692] = `CIPHERTEXT_WIDTH'd4717968;
publickey_row[4693] = `CIPHERTEXT_WIDTH'd16551447;
publickey_row[4694] = `CIPHERTEXT_WIDTH'd6264927;
publickey_row[4695] = `CIPHERTEXT_WIDTH'd6117663;
publickey_row[4696] = `CIPHERTEXT_WIDTH'd9550996;
publickey_row[4697] = `CIPHERTEXT_WIDTH'd5644278;
publickey_row[4698] = `CIPHERTEXT_WIDTH'd4388637;
publickey_row[4699] = `CIPHERTEXT_WIDTH'd2954924;
publickey_row[4700] = `CIPHERTEXT_WIDTH'd12072544;
publickey_row[4701] = `CIPHERTEXT_WIDTH'd8614417;
publickey_row[4702] = `CIPHERTEXT_WIDTH'd12435240;
publickey_row[4703] = `CIPHERTEXT_WIDTH'd3112705;
publickey_row[4704] = `CIPHERTEXT_WIDTH'd11208787;
publickey_row[4705] = `CIPHERTEXT_WIDTH'd11896531;
publickey_row[4706] = `CIPHERTEXT_WIDTH'd1551294;
publickey_row[4707] = `CIPHERTEXT_WIDTH'd4216709;
publickey_row[4708] = `CIPHERTEXT_WIDTH'd1202673;
publickey_row[4709] = `CIPHERTEXT_WIDTH'd10747692;
publickey_row[4710] = `CIPHERTEXT_WIDTH'd1332247;
publickey_row[4711] = `CIPHERTEXT_WIDTH'd14958851;
publickey_row[4712] = `CIPHERTEXT_WIDTH'd14795712;
publickey_row[4713] = `CIPHERTEXT_WIDTH'd3054664;
publickey_row[4714] = `CIPHERTEXT_WIDTH'd16702383;
publickey_row[4715] = `CIPHERTEXT_WIDTH'd9846338;
publickey_row[4716] = `CIPHERTEXT_WIDTH'd10680642;
publickey_row[4717] = `CIPHERTEXT_WIDTH'd6110780;
publickey_row[4718] = `CIPHERTEXT_WIDTH'd7436009;
publickey_row[4719] = `CIPHERTEXT_WIDTH'd4614952;
publickey_row[4720] = `CIPHERTEXT_WIDTH'd18977;
publickey_row[4721] = `CIPHERTEXT_WIDTH'd11836271;
publickey_row[4722] = `CIPHERTEXT_WIDTH'd12636305;
publickey_row[4723] = `CIPHERTEXT_WIDTH'd12768765;
publickey_row[4724] = `CIPHERTEXT_WIDTH'd5613488;
publickey_row[4725] = `CIPHERTEXT_WIDTH'd13788814;
publickey_row[4726] = `CIPHERTEXT_WIDTH'd16224006;
publickey_row[4727] = `CIPHERTEXT_WIDTH'd12556106;
publickey_row[4728] = `CIPHERTEXT_WIDTH'd152666;
publickey_row[4729] = `CIPHERTEXT_WIDTH'd2401279;
publickey_row[4730] = `CIPHERTEXT_WIDTH'd9624319;
publickey_row[4731] = `CIPHERTEXT_WIDTH'd12487518;
publickey_row[4732] = `CIPHERTEXT_WIDTH'd11601360;
publickey_row[4733] = `CIPHERTEXT_WIDTH'd4488933;
publickey_row[4734] = `CIPHERTEXT_WIDTH'd2723258;
publickey_row[4735] = `CIPHERTEXT_WIDTH'd2093275;
publickey_row[4736] = `CIPHERTEXT_WIDTH'd303706;
publickey_row[4737] = `CIPHERTEXT_WIDTH'd399142;
publickey_row[4738] = `CIPHERTEXT_WIDTH'd2350259;
publickey_row[4739] = `CIPHERTEXT_WIDTH'd13420167;
publickey_row[4740] = `CIPHERTEXT_WIDTH'd4871176;
publickey_row[4741] = `CIPHERTEXT_WIDTH'd4603996;
publickey_row[4742] = `CIPHERTEXT_WIDTH'd6705835;
publickey_row[4743] = `CIPHERTEXT_WIDTH'd7812971;
publickey_row[4744] = `CIPHERTEXT_WIDTH'd7502595;
publickey_row[4745] = `CIPHERTEXT_WIDTH'd15152411;
publickey_row[4746] = `CIPHERTEXT_WIDTH'd136793;
publickey_row[4747] = `CIPHERTEXT_WIDTH'd3321482;
publickey_row[4748] = `CIPHERTEXT_WIDTH'd4702470;
publickey_row[4749] = `CIPHERTEXT_WIDTH'd1931587;
publickey_row[4750] = `CIPHERTEXT_WIDTH'd13772438;
publickey_row[4751] = `CIPHERTEXT_WIDTH'd8321227;
publickey_row[4752] = `CIPHERTEXT_WIDTH'd8110741;
publickey_row[4753] = `CIPHERTEXT_WIDTH'd11778722;
publickey_row[4754] = `CIPHERTEXT_WIDTH'd10700204;
publickey_row[4755] = `CIPHERTEXT_WIDTH'd2775296;
publickey_row[4756] = `CIPHERTEXT_WIDTH'd4745284;
publickey_row[4757] = `CIPHERTEXT_WIDTH'd3004658;
publickey_row[4758] = `CIPHERTEXT_WIDTH'd10377651;
publickey_row[4759] = `CIPHERTEXT_WIDTH'd7081574;
publickey_row[4760] = `CIPHERTEXT_WIDTH'd15217206;
publickey_row[4761] = `CIPHERTEXT_WIDTH'd7027435;
publickey_row[4762] = `CIPHERTEXT_WIDTH'd4643829;
publickey_row[4763] = `CIPHERTEXT_WIDTH'd11305469;
publickey_row[4764] = `CIPHERTEXT_WIDTH'd15008070;
publickey_row[4765] = `CIPHERTEXT_WIDTH'd12979320;
publickey_row[4766] = `CIPHERTEXT_WIDTH'd7198777;
publickey_row[4767] = `CIPHERTEXT_WIDTH'd12115384;
publickey_row[4768] = `CIPHERTEXT_WIDTH'd8578252;
publickey_row[4769] = `CIPHERTEXT_WIDTH'd9324792;
publickey_row[4770] = `CIPHERTEXT_WIDTH'd5245197;
publickey_row[4771] = `CIPHERTEXT_WIDTH'd15349223;
publickey_row[4772] = `CIPHERTEXT_WIDTH'd7726059;
publickey_row[4773] = `CIPHERTEXT_WIDTH'd13964207;
publickey_row[4774] = `CIPHERTEXT_WIDTH'd345620;
publickey_row[4775] = `CIPHERTEXT_WIDTH'd8584751;
publickey_row[4776] = `CIPHERTEXT_WIDTH'd13762763;
publickey_row[4777] = `CIPHERTEXT_WIDTH'd2617649;
publickey_row[4778] = `CIPHERTEXT_WIDTH'd14728537;
publickey_row[4779] = `CIPHERTEXT_WIDTH'd9491940;
publickey_row[4780] = `CIPHERTEXT_WIDTH'd4184925;
publickey_row[4781] = `CIPHERTEXT_WIDTH'd13595522;
publickey_row[4782] = `CIPHERTEXT_WIDTH'd658539;
publickey_row[4783] = `CIPHERTEXT_WIDTH'd8525426;
publickey_row[4784] = `CIPHERTEXT_WIDTH'd53063;
publickey_row[4785] = `CIPHERTEXT_WIDTH'd5050351;
publickey_row[4786] = `CIPHERTEXT_WIDTH'd2618679;
publickey_row[4787] = `CIPHERTEXT_WIDTH'd2144911;
publickey_row[4788] = `CIPHERTEXT_WIDTH'd7589545;
publickey_row[4789] = `CIPHERTEXT_WIDTH'd3661080;
publickey_row[4790] = `CIPHERTEXT_WIDTH'd5421013;
publickey_row[4791] = `CIPHERTEXT_WIDTH'd11881040;
publickey_row[4792] = `CIPHERTEXT_WIDTH'd5219227;
publickey_row[4793] = `CIPHERTEXT_WIDTH'd4187332;
publickey_row[4794] = `CIPHERTEXT_WIDTH'd6694213;
publickey_row[4795] = `CIPHERTEXT_WIDTH'd12369494;
publickey_row[4796] = `CIPHERTEXT_WIDTH'd8766895;
publickey_row[4797] = `CIPHERTEXT_WIDTH'd4340089;
publickey_row[4798] = `CIPHERTEXT_WIDTH'd11959058;
publickey_row[4799] = `CIPHERTEXT_WIDTH'd13218674;
publickey_row[4800] = `CIPHERTEXT_WIDTH'd4842431;
publickey_row[4801] = `CIPHERTEXT_WIDTH'd10827724;
publickey_row[4802] = `CIPHERTEXT_WIDTH'd11600617;
publickey_row[4803] = `CIPHERTEXT_WIDTH'd4088436;
publickey_row[4804] = `CIPHERTEXT_WIDTH'd1900454;
publickey_row[4805] = `CIPHERTEXT_WIDTH'd5225855;
publickey_row[4806] = `CIPHERTEXT_WIDTH'd10291726;
publickey_row[4807] = `CIPHERTEXT_WIDTH'd4394865;
publickey_row[4808] = `CIPHERTEXT_WIDTH'd5067562;
publickey_row[4809] = `CIPHERTEXT_WIDTH'd9101257;
publickey_row[4810] = `CIPHERTEXT_WIDTH'd627699;
publickey_row[4811] = `CIPHERTEXT_WIDTH'd11462657;
publickey_row[4812] = `CIPHERTEXT_WIDTH'd12392880;
publickey_row[4813] = `CIPHERTEXT_WIDTH'd7579656;
publickey_row[4814] = `CIPHERTEXT_WIDTH'd204034;
publickey_row[4815] = `CIPHERTEXT_WIDTH'd5278471;
publickey_row[4816] = `CIPHERTEXT_WIDTH'd15117340;
publickey_row[4817] = `CIPHERTEXT_WIDTH'd9845724;
publickey_row[4818] = `CIPHERTEXT_WIDTH'd12812714;
publickey_row[4819] = `CIPHERTEXT_WIDTH'd3583249;
publickey_row[4820] = `CIPHERTEXT_WIDTH'd2698238;
publickey_row[4821] = `CIPHERTEXT_WIDTH'd12918609;
publickey_row[4822] = `CIPHERTEXT_WIDTH'd13085686;
publickey_row[4823] = `CIPHERTEXT_WIDTH'd13551044;
publickey_row[4824] = `CIPHERTEXT_WIDTH'd5749961;
publickey_row[4825] = `CIPHERTEXT_WIDTH'd3065205;
publickey_row[4826] = `CIPHERTEXT_WIDTH'd5594481;
publickey_row[4827] = `CIPHERTEXT_WIDTH'd8877377;
publickey_row[4828] = `CIPHERTEXT_WIDTH'd5548095;
publickey_row[4829] = `CIPHERTEXT_WIDTH'd15413164;
publickey_row[4830] = `CIPHERTEXT_WIDTH'd10641144;
publickey_row[4831] = `CIPHERTEXT_WIDTH'd3609839;
publickey_row[4832] = `CIPHERTEXT_WIDTH'd12719580;
publickey_row[4833] = `CIPHERTEXT_WIDTH'd9998474;
publickey_row[4834] = `CIPHERTEXT_WIDTH'd1747534;
publickey_row[4835] = `CIPHERTEXT_WIDTH'd3545900;
publickey_row[4836] = `CIPHERTEXT_WIDTH'd15057909;
publickey_row[4837] = `CIPHERTEXT_WIDTH'd14893381;
publickey_row[4838] = `CIPHERTEXT_WIDTH'd13012793;
publickey_row[4839] = `CIPHERTEXT_WIDTH'd8100588;
publickey_row[4840] = `CIPHERTEXT_WIDTH'd9068024;
publickey_row[4841] = `CIPHERTEXT_WIDTH'd8390695;
publickey_row[4842] = `CIPHERTEXT_WIDTH'd7516557;
publickey_row[4843] = `CIPHERTEXT_WIDTH'd12087689;
publickey_row[4844] = `CIPHERTEXT_WIDTH'd2356042;
publickey_row[4845] = `CIPHERTEXT_WIDTH'd13439114;
publickey_row[4846] = `CIPHERTEXT_WIDTH'd6045557;
publickey_row[4847] = `CIPHERTEXT_WIDTH'd3619051;
publickey_row[4848] = `CIPHERTEXT_WIDTH'd4968884;
publickey_row[4849] = `CIPHERTEXT_WIDTH'd5283595;
publickey_row[4850] = `CIPHERTEXT_WIDTH'd6181151;
publickey_row[4851] = `CIPHERTEXT_WIDTH'd15348582;
publickey_row[4852] = `CIPHERTEXT_WIDTH'd12725641;
publickey_row[4853] = `CIPHERTEXT_WIDTH'd11245223;
publickey_row[4854] = `CIPHERTEXT_WIDTH'd12661408;
publickey_row[4855] = `CIPHERTEXT_WIDTH'd16706004;
publickey_row[4856] = `CIPHERTEXT_WIDTH'd13276763;
publickey_row[4857] = `CIPHERTEXT_WIDTH'd1660046;
publickey_row[4858] = `CIPHERTEXT_WIDTH'd16670492;
publickey_row[4859] = `CIPHERTEXT_WIDTH'd2352891;
publickey_row[4860] = `CIPHERTEXT_WIDTH'd10877672;
publickey_row[4861] = `CIPHERTEXT_WIDTH'd9460852;
publickey_row[4862] = `CIPHERTEXT_WIDTH'd847477;
publickey_row[4863] = `CIPHERTEXT_WIDTH'd12821964;
publickey_row[4864] = `CIPHERTEXT_WIDTH'd1687463;
publickey_row[4865] = `CIPHERTEXT_WIDTH'd14917744;
publickey_row[4866] = `CIPHERTEXT_WIDTH'd13035204;
publickey_row[4867] = `CIPHERTEXT_WIDTH'd15674661;
publickey_row[4868] = `CIPHERTEXT_WIDTH'd12840916;
publickey_row[4869] = `CIPHERTEXT_WIDTH'd4975518;
publickey_row[4870] = `CIPHERTEXT_WIDTH'd4899136;
publickey_row[4871] = `CIPHERTEXT_WIDTH'd14262911;
publickey_row[4872] = `CIPHERTEXT_WIDTH'd14605285;
publickey_row[4873] = `CIPHERTEXT_WIDTH'd554568;
publickey_row[4874] = `CIPHERTEXT_WIDTH'd1295217;
publickey_row[4875] = `CIPHERTEXT_WIDTH'd1391800;
publickey_row[4876] = `CIPHERTEXT_WIDTH'd732233;
publickey_row[4877] = `CIPHERTEXT_WIDTH'd5752692;
publickey_row[4878] = `CIPHERTEXT_WIDTH'd4902241;
publickey_row[4879] = `CIPHERTEXT_WIDTH'd4610834;
publickey_row[4880] = `CIPHERTEXT_WIDTH'd4598123;
publickey_row[4881] = `CIPHERTEXT_WIDTH'd9185652;
publickey_row[4882] = `CIPHERTEXT_WIDTH'd5305552;
publickey_row[4883] = `CIPHERTEXT_WIDTH'd6341304;
publickey_row[4884] = `CIPHERTEXT_WIDTH'd10376122;
publickey_row[4885] = `CIPHERTEXT_WIDTH'd11282637;
publickey_row[4886] = `CIPHERTEXT_WIDTH'd9922194;
publickey_row[4887] = `CIPHERTEXT_WIDTH'd10433922;
publickey_row[4888] = `CIPHERTEXT_WIDTH'd12548277;
publickey_row[4889] = `CIPHERTEXT_WIDTH'd7128142;
publickey_row[4890] = `CIPHERTEXT_WIDTH'd6648039;
publickey_row[4891] = `CIPHERTEXT_WIDTH'd5054205;
publickey_row[4892] = `CIPHERTEXT_WIDTH'd4451173;
publickey_row[4893] = `CIPHERTEXT_WIDTH'd3922665;
publickey_row[4894] = `CIPHERTEXT_WIDTH'd10799385;
publickey_row[4895] = `CIPHERTEXT_WIDTH'd2934044;
publickey_row[4896] = `CIPHERTEXT_WIDTH'd11277752;
publickey_row[4897] = `CIPHERTEXT_WIDTH'd5413420;
publickey_row[4898] = `CIPHERTEXT_WIDTH'd9821733;
publickey_row[4899] = `CIPHERTEXT_WIDTH'd3116509;
publickey_row[4900] = `CIPHERTEXT_WIDTH'd10083521;
publickey_row[4901] = `CIPHERTEXT_WIDTH'd12976393;
publickey_row[4902] = `CIPHERTEXT_WIDTH'd1844279;
publickey_row[4903] = `CIPHERTEXT_WIDTH'd997852;
publickey_row[4904] = `CIPHERTEXT_WIDTH'd1738362;
publickey_row[4905] = `CIPHERTEXT_WIDTH'd4924420;
publickey_row[4906] = `CIPHERTEXT_WIDTH'd9085437;
publickey_row[4907] = `CIPHERTEXT_WIDTH'd15241316;
publickey_row[4908] = `CIPHERTEXT_WIDTH'd5194195;
publickey_row[4909] = `CIPHERTEXT_WIDTH'd16445496;
publickey_row[4910] = `CIPHERTEXT_WIDTH'd2729138;
publickey_row[4911] = `CIPHERTEXT_WIDTH'd5317736;
publickey_row[4912] = `CIPHERTEXT_WIDTH'd5401397;
publickey_row[4913] = `CIPHERTEXT_WIDTH'd8833374;
publickey_row[4914] = `CIPHERTEXT_WIDTH'd964165;
publickey_row[4915] = `CIPHERTEXT_WIDTH'd4141494;
publickey_row[4916] = `CIPHERTEXT_WIDTH'd10882298;
publickey_row[4917] = `CIPHERTEXT_WIDTH'd5773341;
publickey_row[4918] = `CIPHERTEXT_WIDTH'd9674206;
publickey_row[4919] = `CIPHERTEXT_WIDTH'd1999483;
publickey_row[4920] = `CIPHERTEXT_WIDTH'd9652571;
publickey_row[4921] = `CIPHERTEXT_WIDTH'd4776231;
publickey_row[4922] = `CIPHERTEXT_WIDTH'd5561126;
publickey_row[4923] = `CIPHERTEXT_WIDTH'd3274444;
publickey_row[4924] = `CIPHERTEXT_WIDTH'd8157225;
publickey_row[4925] = `CIPHERTEXT_WIDTH'd12089227;
publickey_row[4926] = `CIPHERTEXT_WIDTH'd9224515;
publickey_row[4927] = `CIPHERTEXT_WIDTH'd5191397;
publickey_row[4928] = `CIPHERTEXT_WIDTH'd2261099;
publickey_row[4929] = `CIPHERTEXT_WIDTH'd5907304;
publickey_row[4930] = `CIPHERTEXT_WIDTH'd2890162;
publickey_row[4931] = `CIPHERTEXT_WIDTH'd7962516;
publickey_row[4932] = `CIPHERTEXT_WIDTH'd10337304;
publickey_row[4933] = `CIPHERTEXT_WIDTH'd5179911;
publickey_row[4934] = `CIPHERTEXT_WIDTH'd1135251;
publickey_row[4935] = `CIPHERTEXT_WIDTH'd10964503;
publickey_row[4936] = `CIPHERTEXT_WIDTH'd12911154;
publickey_row[4937] = `CIPHERTEXT_WIDTH'd15690726;
publickey_row[4938] = `CIPHERTEXT_WIDTH'd15571940;
publickey_row[4939] = `CIPHERTEXT_WIDTH'd2069229;
publickey_row[4940] = `CIPHERTEXT_WIDTH'd5047981;
publickey_row[4941] = `CIPHERTEXT_WIDTH'd7174039;
publickey_row[4942] = `CIPHERTEXT_WIDTH'd4894755;
publickey_row[4943] = `CIPHERTEXT_WIDTH'd781113;
publickey_row[4944] = `CIPHERTEXT_WIDTH'd10468667;
publickey_row[4945] = `CIPHERTEXT_WIDTH'd7896696;
publickey_row[4946] = `CIPHERTEXT_WIDTH'd4641139;
publickey_row[4947] = `CIPHERTEXT_WIDTH'd5698724;
publickey_row[4948] = `CIPHERTEXT_WIDTH'd12499842;
publickey_row[4949] = `CIPHERTEXT_WIDTH'd15712920;
publickey_row[4950] = `CIPHERTEXT_WIDTH'd4428658;
publickey_row[4951] = `CIPHERTEXT_WIDTH'd12831895;
publickey_row[4952] = `CIPHERTEXT_WIDTH'd8253340;
publickey_row[4953] = `CIPHERTEXT_WIDTH'd14227470;
publickey_row[4954] = `CIPHERTEXT_WIDTH'd8070239;
publickey_row[4955] = `CIPHERTEXT_WIDTH'd15615812;
publickey_row[4956] = `CIPHERTEXT_WIDTH'd12042975;
publickey_row[4957] = `CIPHERTEXT_WIDTH'd2965798;
publickey_row[4958] = `CIPHERTEXT_WIDTH'd7508620;
publickey_row[4959] = `CIPHERTEXT_WIDTH'd15076929;
publickey_row[4960] = `CIPHERTEXT_WIDTH'd1080646;
publickey_row[4961] = `CIPHERTEXT_WIDTH'd5681103;
publickey_row[4962] = `CIPHERTEXT_WIDTH'd381587;
publickey_row[4963] = `CIPHERTEXT_WIDTH'd10759280;
publickey_row[4964] = `CIPHERTEXT_WIDTH'd16328469;
publickey_row[4965] = `CIPHERTEXT_WIDTH'd165972;
publickey_row[4966] = `CIPHERTEXT_WIDTH'd8813108;
publickey_row[4967] = `CIPHERTEXT_WIDTH'd109390;
publickey_row[4968] = `CIPHERTEXT_WIDTH'd16176175;
publickey_row[4969] = `CIPHERTEXT_WIDTH'd13382782;
publickey_row[4970] = `CIPHERTEXT_WIDTH'd5587287;
publickey_row[4971] = `CIPHERTEXT_WIDTH'd13313268;
publickey_row[4972] = `CIPHERTEXT_WIDTH'd2020572;
publickey_row[4973] = `CIPHERTEXT_WIDTH'd1661280;
publickey_row[4974] = `CIPHERTEXT_WIDTH'd2929554;
publickey_row[4975] = `CIPHERTEXT_WIDTH'd8474521;
publickey_row[4976] = `CIPHERTEXT_WIDTH'd8245340;
publickey_row[4977] = `CIPHERTEXT_WIDTH'd1517601;
publickey_row[4978] = `CIPHERTEXT_WIDTH'd13106588;
publickey_row[4979] = `CIPHERTEXT_WIDTH'd13856160;
publickey_row[4980] = `CIPHERTEXT_WIDTH'd3702189;
publickey_row[4981] = `CIPHERTEXT_WIDTH'd6864036;
publickey_row[4982] = `CIPHERTEXT_WIDTH'd15986398;
publickey_row[4983] = `CIPHERTEXT_WIDTH'd7555844;
publickey_row[4984] = `CIPHERTEXT_WIDTH'd9001661;
publickey_row[4985] = `CIPHERTEXT_WIDTH'd14359306;
publickey_row[4986] = `CIPHERTEXT_WIDTH'd2284291;
publickey_row[4987] = `CIPHERTEXT_WIDTH'd11723153;
publickey_row[4988] = `CIPHERTEXT_WIDTH'd5672208;
publickey_row[4989] = `CIPHERTEXT_WIDTH'd3064186;
publickey_row[4990] = `CIPHERTEXT_WIDTH'd8263459;
publickey_row[4991] = `CIPHERTEXT_WIDTH'd7637725;
publickey_row[4992] = `CIPHERTEXT_WIDTH'd11219425;
publickey_row[4993] = `CIPHERTEXT_WIDTH'd12717002;
publickey_row[4994] = `CIPHERTEXT_WIDTH'd7065732;
publickey_row[4995] = `CIPHERTEXT_WIDTH'd16201930;
publickey_row[4996] = `CIPHERTEXT_WIDTH'd3706442;
publickey_row[4997] = `CIPHERTEXT_WIDTH'd5324855;
publickey_row[4998] = `CIPHERTEXT_WIDTH'd5327117;
publickey_row[4999] = `CIPHERTEXT_WIDTH'd13290099;
publickey_row[5000] = `CIPHERTEXT_WIDTH'd9423544;
publickey_row[5001] = `CIPHERTEXT_WIDTH'd7385945;
publickey_row[5002] = `CIPHERTEXT_WIDTH'd6387033;
publickey_row[5003] = `CIPHERTEXT_WIDTH'd2029569;
publickey_row[5004] = `CIPHERTEXT_WIDTH'd10579921;
publickey_row[5005] = `CIPHERTEXT_WIDTH'd4068161;
publickey_row[5006] = `CIPHERTEXT_WIDTH'd14551;
publickey_row[5007] = `CIPHERTEXT_WIDTH'd16339133;
publickey_row[5008] = `CIPHERTEXT_WIDTH'd10467803;
publickey_row[5009] = `CIPHERTEXT_WIDTH'd5671163;
publickey_row[5010] = `CIPHERTEXT_WIDTH'd12404238;
publickey_row[5011] = `CIPHERTEXT_WIDTH'd4900622;
publickey_row[5012] = `CIPHERTEXT_WIDTH'd8332782;
publickey_row[5013] = `CIPHERTEXT_WIDTH'd14321202;
publickey_row[5014] = `CIPHERTEXT_WIDTH'd11361664;
publickey_row[5015] = `CIPHERTEXT_WIDTH'd11335357;
publickey_row[5016] = `CIPHERTEXT_WIDTH'd7284058;
publickey_row[5017] = `CIPHERTEXT_WIDTH'd11581784;
publickey_row[5018] = `CIPHERTEXT_WIDTH'd6378173;
publickey_row[5019] = `CIPHERTEXT_WIDTH'd13954894;
publickey_row[5020] = `CIPHERTEXT_WIDTH'd6493226;
publickey_row[5021] = `CIPHERTEXT_WIDTH'd8354300;
publickey_row[5022] = `CIPHERTEXT_WIDTH'd11780614;
publickey_row[5023] = `CIPHERTEXT_WIDTH'd9428926;
publickey_row[5024] = `CIPHERTEXT_WIDTH'd4208386;
publickey_row[5025] = `CIPHERTEXT_WIDTH'd9538025;
publickey_row[5026] = `CIPHERTEXT_WIDTH'd13342548;
publickey_row[5027] = `CIPHERTEXT_WIDTH'd661445;
publickey_row[5028] = `CIPHERTEXT_WIDTH'd7831527;
publickey_row[5029] = `CIPHERTEXT_WIDTH'd11192119;
publickey_row[5030] = `CIPHERTEXT_WIDTH'd4168315;
publickey_row[5031] = `CIPHERTEXT_WIDTH'd5124508;
publickey_row[5032] = `CIPHERTEXT_WIDTH'd19425;
publickey_row[5033] = `CIPHERTEXT_WIDTH'd13344221;
publickey_row[5034] = `CIPHERTEXT_WIDTH'd2680548;
publickey_row[5035] = `CIPHERTEXT_WIDTH'd14347403;
publickey_row[5036] = `CIPHERTEXT_WIDTH'd2890294;
publickey_row[5037] = `CIPHERTEXT_WIDTH'd10234197;
publickey_row[5038] = `CIPHERTEXT_WIDTH'd11796751;
publickey_row[5039] = `CIPHERTEXT_WIDTH'd4918976;
publickey_row[5040] = `CIPHERTEXT_WIDTH'd6523501;
publickey_row[5041] = `CIPHERTEXT_WIDTH'd4903167;
publickey_row[5042] = `CIPHERTEXT_WIDTH'd1499816;
publickey_row[5043] = `CIPHERTEXT_WIDTH'd5197468;
publickey_row[5044] = `CIPHERTEXT_WIDTH'd3514389;
publickey_row[5045] = `CIPHERTEXT_WIDTH'd12318019;
publickey_row[5046] = `CIPHERTEXT_WIDTH'd8549479;
publickey_row[5047] = `CIPHERTEXT_WIDTH'd5334366;
publickey_row[5048] = `CIPHERTEXT_WIDTH'd15643310;
publickey_row[5049] = `CIPHERTEXT_WIDTH'd7762975;
publickey_row[5050] = `CIPHERTEXT_WIDTH'd4993057;
publickey_row[5051] = `CIPHERTEXT_WIDTH'd13371024;
publickey_row[5052] = `CIPHERTEXT_WIDTH'd8471425;
publickey_row[5053] = `CIPHERTEXT_WIDTH'd10943338;
publickey_row[5054] = `CIPHERTEXT_WIDTH'd11880113;
publickey_row[5055] = `CIPHERTEXT_WIDTH'd1801830;
publickey_row[5056] = `CIPHERTEXT_WIDTH'd8340364;
publickey_row[5057] = `CIPHERTEXT_WIDTH'd8886277;
publickey_row[5058] = `CIPHERTEXT_WIDTH'd255555;
publickey_row[5059] = `CIPHERTEXT_WIDTH'd9743181;
publickey_row[5060] = `CIPHERTEXT_WIDTH'd9474011;
publickey_row[5061] = `CIPHERTEXT_WIDTH'd7584215;
publickey_row[5062] = `CIPHERTEXT_WIDTH'd2721472;
publickey_row[5063] = `CIPHERTEXT_WIDTH'd13093938;
publickey_row[5064] = `CIPHERTEXT_WIDTH'd841704;
publickey_row[5065] = `CIPHERTEXT_WIDTH'd2681614;
publickey_row[5066] = `CIPHERTEXT_WIDTH'd210066;
publickey_row[5067] = `CIPHERTEXT_WIDTH'd12347030;
publickey_row[5068] = `CIPHERTEXT_WIDTH'd7219972;
publickey_row[5069] = `CIPHERTEXT_WIDTH'd11543063;
publickey_row[5070] = `CIPHERTEXT_WIDTH'd15617439;
publickey_row[5071] = `CIPHERTEXT_WIDTH'd3360431;
publickey_row[5072] = `CIPHERTEXT_WIDTH'd698175;
publickey_row[5073] = `CIPHERTEXT_WIDTH'd388018;
publickey_row[5074] = `CIPHERTEXT_WIDTH'd4277838;
publickey_row[5075] = `CIPHERTEXT_WIDTH'd4687107;
publickey_row[5076] = `CIPHERTEXT_WIDTH'd14279331;
publickey_row[5077] = `CIPHERTEXT_WIDTH'd4841122;
publickey_row[5078] = `CIPHERTEXT_WIDTH'd15219834;
publickey_row[5079] = `CIPHERTEXT_WIDTH'd15032604;
publickey_row[5080] = `CIPHERTEXT_WIDTH'd1224306;
publickey_row[5081] = `CIPHERTEXT_WIDTH'd9734647;
publickey_row[5082] = `CIPHERTEXT_WIDTH'd8759539;
publickey_row[5083] = `CIPHERTEXT_WIDTH'd14137287;
publickey_row[5084] = `CIPHERTEXT_WIDTH'd9883659;
publickey_row[5085] = `CIPHERTEXT_WIDTH'd7018954;
publickey_row[5086] = `CIPHERTEXT_WIDTH'd3549312;
publickey_row[5087] = `CIPHERTEXT_WIDTH'd4573056;
publickey_row[5088] = `CIPHERTEXT_WIDTH'd6463186;
publickey_row[5089] = `CIPHERTEXT_WIDTH'd14536015;
publickey_row[5090] = `CIPHERTEXT_WIDTH'd31118;
publickey_row[5091] = `CIPHERTEXT_WIDTH'd16073486;
publickey_row[5092] = `CIPHERTEXT_WIDTH'd11028103;
publickey_row[5093] = `CIPHERTEXT_WIDTH'd12708885;
publickey_row[5094] = `CIPHERTEXT_WIDTH'd13625560;
publickey_row[5095] = `CIPHERTEXT_WIDTH'd11990846;
publickey_row[5096] = `CIPHERTEXT_WIDTH'd12272993;
publickey_row[5097] = `CIPHERTEXT_WIDTH'd1488881;
publickey_row[5098] = `CIPHERTEXT_WIDTH'd12090340;
publickey_row[5099] = `CIPHERTEXT_WIDTH'd14013607;
publickey_row[5100] = `CIPHERTEXT_WIDTH'd3872611;
publickey_row[5101] = `CIPHERTEXT_WIDTH'd10926032;
publickey_row[5102] = `CIPHERTEXT_WIDTH'd9830228;
publickey_row[5103] = `CIPHERTEXT_WIDTH'd2889379;
publickey_row[5104] = `CIPHERTEXT_WIDTH'd6322728;
publickey_row[5105] = `CIPHERTEXT_WIDTH'd10503119;
publickey_row[5106] = `CIPHERTEXT_WIDTH'd14935143;
publickey_row[5107] = `CIPHERTEXT_WIDTH'd9169177;
publickey_row[5108] = `CIPHERTEXT_WIDTH'd4195671;
publickey_row[5109] = `CIPHERTEXT_WIDTH'd1675930;
publickey_row[5110] = `CIPHERTEXT_WIDTH'd13139693;
publickey_row[5111] = `CIPHERTEXT_WIDTH'd4801989;
publickey_row[5112] = `CIPHERTEXT_WIDTH'd14631537;
publickey_row[5113] = `CIPHERTEXT_WIDTH'd13671528;
publickey_row[5114] = `CIPHERTEXT_WIDTH'd12902088;
publickey_row[5115] = `CIPHERTEXT_WIDTH'd4610827;
publickey_row[5116] = `CIPHERTEXT_WIDTH'd16515004;
publickey_row[5117] = `CIPHERTEXT_WIDTH'd246446;
publickey_row[5118] = `CIPHERTEXT_WIDTH'd611867;
publickey_row[5119] = `CIPHERTEXT_WIDTH'd3154240;
publickey_row[5120] = `CIPHERTEXT_WIDTH'd8572628;
publickey_row[5121] = `CIPHERTEXT_WIDTH'd2184393;
publickey_row[5122] = `CIPHERTEXT_WIDTH'd12786536;
publickey_row[5123] = `CIPHERTEXT_WIDTH'd7415072;
publickey_row[5124] = `CIPHERTEXT_WIDTH'd10488761;
publickey_row[5125] = `CIPHERTEXT_WIDTH'd7049550;
publickey_row[5126] = `CIPHERTEXT_WIDTH'd1399861;
publickey_row[5127] = `CIPHERTEXT_WIDTH'd2681548;
publickey_row[5128] = `CIPHERTEXT_WIDTH'd8950263;
publickey_row[5129] = `CIPHERTEXT_WIDTH'd327054;
publickey_row[5130] = `CIPHERTEXT_WIDTH'd7557845;
publickey_row[5131] = `CIPHERTEXT_WIDTH'd15598863;
publickey_row[5132] = `CIPHERTEXT_WIDTH'd13801121;
publickey_row[5133] = `CIPHERTEXT_WIDTH'd4622050;
publickey_row[5134] = `CIPHERTEXT_WIDTH'd748981;
publickey_row[5135] = `CIPHERTEXT_WIDTH'd16557353;
publickey_row[5136] = `CIPHERTEXT_WIDTH'd11476680;
publickey_row[5137] = `CIPHERTEXT_WIDTH'd10841563;
publickey_row[5138] = `CIPHERTEXT_WIDTH'd11219211;
publickey_row[5139] = `CIPHERTEXT_WIDTH'd14240137;
publickey_row[5140] = `CIPHERTEXT_WIDTH'd13654239;
publickey_row[5141] = `CIPHERTEXT_WIDTH'd10298731;
publickey_row[5142] = `CIPHERTEXT_WIDTH'd237466;
publickey_row[5143] = `CIPHERTEXT_WIDTH'd1854644;
publickey_row[5144] = `CIPHERTEXT_WIDTH'd2930741;
publickey_row[5145] = `CIPHERTEXT_WIDTH'd12275199;
publickey_row[5146] = `CIPHERTEXT_WIDTH'd11640205;
publickey_row[5147] = `CIPHERTEXT_WIDTH'd15162122;
publickey_row[5148] = `CIPHERTEXT_WIDTH'd2536720;
publickey_row[5149] = `CIPHERTEXT_WIDTH'd2874053;
publickey_row[5150] = `CIPHERTEXT_WIDTH'd3480546;
publickey_row[5151] = `CIPHERTEXT_WIDTH'd2665766;
publickey_row[5152] = `CIPHERTEXT_WIDTH'd80148;
publickey_row[5153] = `CIPHERTEXT_WIDTH'd1605472;
publickey_row[5154] = `CIPHERTEXT_WIDTH'd4864668;
publickey_row[5155] = `CIPHERTEXT_WIDTH'd16262984;
publickey_row[5156] = `CIPHERTEXT_WIDTH'd12943506;
publickey_row[5157] = `CIPHERTEXT_WIDTH'd943509;
publickey_row[5158] = `CIPHERTEXT_WIDTH'd7615614;
publickey_row[5159] = `CIPHERTEXT_WIDTH'd1614867;
publickey_row[5160] = `CIPHERTEXT_WIDTH'd7348079;
publickey_row[5161] = `CIPHERTEXT_WIDTH'd3164233;
publickey_row[5162] = `CIPHERTEXT_WIDTH'd6287672;
publickey_row[5163] = `CIPHERTEXT_WIDTH'd2302670;
publickey_row[5164] = `CIPHERTEXT_WIDTH'd6134111;
publickey_row[5165] = `CIPHERTEXT_WIDTH'd8072049;
publickey_row[5166] = `CIPHERTEXT_WIDTH'd13238839;
publickey_row[5167] = `CIPHERTEXT_WIDTH'd7321885;
publickey_row[5168] = `CIPHERTEXT_WIDTH'd6424659;
publickey_row[5169] = `CIPHERTEXT_WIDTH'd16379596;
publickey_row[5170] = `CIPHERTEXT_WIDTH'd2763569;
publickey_row[5171] = `CIPHERTEXT_WIDTH'd5787913;
publickey_row[5172] = `CIPHERTEXT_WIDTH'd15404759;
publickey_row[5173] = `CIPHERTEXT_WIDTH'd3507625;
publickey_row[5174] = `CIPHERTEXT_WIDTH'd5918651;
publickey_row[5175] = `CIPHERTEXT_WIDTH'd8208175;
publickey_row[5176] = `CIPHERTEXT_WIDTH'd7473130;
publickey_row[5177] = `CIPHERTEXT_WIDTH'd13238147;
publickey_row[5178] = `CIPHERTEXT_WIDTH'd649391;
publickey_row[5179] = `CIPHERTEXT_WIDTH'd16338078;
publickey_row[5180] = `CIPHERTEXT_WIDTH'd15896656;
publickey_row[5181] = `CIPHERTEXT_WIDTH'd2187953;
publickey_row[5182] = `CIPHERTEXT_WIDTH'd9020310;
publickey_row[5183] = `CIPHERTEXT_WIDTH'd5441572;
publickey_row[5184] = `CIPHERTEXT_WIDTH'd10058693;
publickey_row[5185] = `CIPHERTEXT_WIDTH'd2687874;
publickey_row[5186] = `CIPHERTEXT_WIDTH'd13468299;
publickey_row[5187] = `CIPHERTEXT_WIDTH'd8034673;
publickey_row[5188] = `CIPHERTEXT_WIDTH'd6824920;
publickey_row[5189] = `CIPHERTEXT_WIDTH'd7444137;
publickey_row[5190] = `CIPHERTEXT_WIDTH'd16268905;
publickey_row[5191] = `CIPHERTEXT_WIDTH'd15533998;
publickey_row[5192] = `CIPHERTEXT_WIDTH'd5272764;
publickey_row[5193] = `CIPHERTEXT_WIDTH'd12409978;
publickey_row[5194] = `CIPHERTEXT_WIDTH'd9268006;
publickey_row[5195] = `CIPHERTEXT_WIDTH'd16338523;
publickey_row[5196] = `CIPHERTEXT_WIDTH'd3623389;
publickey_row[5197] = `CIPHERTEXT_WIDTH'd5956883;
publickey_row[5198] = `CIPHERTEXT_WIDTH'd16346131;
publickey_row[5199] = `CIPHERTEXT_WIDTH'd7119480;
publickey_row[5200] = `CIPHERTEXT_WIDTH'd1585308;
publickey_row[5201] = `CIPHERTEXT_WIDTH'd2173243;
publickey_row[5202] = `CIPHERTEXT_WIDTH'd724143;
publickey_row[5203] = `CIPHERTEXT_WIDTH'd4945326;
publickey_row[5204] = `CIPHERTEXT_WIDTH'd6815089;
publickey_row[5205] = `CIPHERTEXT_WIDTH'd8762555;
publickey_row[5206] = `CIPHERTEXT_WIDTH'd2489518;
publickey_row[5207] = `CIPHERTEXT_WIDTH'd16280329;
publickey_row[5208] = `CIPHERTEXT_WIDTH'd15359391;
publickey_row[5209] = `CIPHERTEXT_WIDTH'd3014882;
publickey_row[5210] = `CIPHERTEXT_WIDTH'd6991161;
publickey_row[5211] = `CIPHERTEXT_WIDTH'd6327606;
publickey_row[5212] = `CIPHERTEXT_WIDTH'd2469136;
publickey_row[5213] = `CIPHERTEXT_WIDTH'd3852408;
publickey_row[5214] = `CIPHERTEXT_WIDTH'd3180935;
publickey_row[5215] = `CIPHERTEXT_WIDTH'd5964341;
publickey_row[5216] = `CIPHERTEXT_WIDTH'd11362986;
publickey_row[5217] = `CIPHERTEXT_WIDTH'd4749137;
publickey_row[5218] = `CIPHERTEXT_WIDTH'd5149952;
publickey_row[5219] = `CIPHERTEXT_WIDTH'd8596740;
publickey_row[5220] = `CIPHERTEXT_WIDTH'd4428147;
publickey_row[5221] = `CIPHERTEXT_WIDTH'd2285398;
publickey_row[5222] = `CIPHERTEXT_WIDTH'd8136405;
publickey_row[5223] = `CIPHERTEXT_WIDTH'd9801447;
publickey_row[5224] = `CIPHERTEXT_WIDTH'd468957;
publickey_row[5225] = `CIPHERTEXT_WIDTH'd14672412;
publickey_row[5226] = `CIPHERTEXT_WIDTH'd5984890;
publickey_row[5227] = `CIPHERTEXT_WIDTH'd10871466;
publickey_row[5228] = `CIPHERTEXT_WIDTH'd1912391;
publickey_row[5229] = `CIPHERTEXT_WIDTH'd6550025;
publickey_row[5230] = `CIPHERTEXT_WIDTH'd12023543;
publickey_row[5231] = `CIPHERTEXT_WIDTH'd6155473;
publickey_row[5232] = `CIPHERTEXT_WIDTH'd7932029;
publickey_row[5233] = `CIPHERTEXT_WIDTH'd613116;
publickey_row[5234] = `CIPHERTEXT_WIDTH'd14147759;
publickey_row[5235] = `CIPHERTEXT_WIDTH'd4488251;
publickey_row[5236] = `CIPHERTEXT_WIDTH'd6967062;
publickey_row[5237] = `CIPHERTEXT_WIDTH'd9616470;
publickey_row[5238] = `CIPHERTEXT_WIDTH'd10876032;
publickey_row[5239] = `CIPHERTEXT_WIDTH'd11936682;
publickey_row[5240] = `CIPHERTEXT_WIDTH'd9431329;
publickey_row[5241] = `CIPHERTEXT_WIDTH'd16491081;
publickey_row[5242] = `CIPHERTEXT_WIDTH'd8627797;
publickey_row[5243] = `CIPHERTEXT_WIDTH'd15333159;
publickey_row[5244] = `CIPHERTEXT_WIDTH'd278733;
publickey_row[5245] = `CIPHERTEXT_WIDTH'd11270891;
publickey_row[5246] = `CIPHERTEXT_WIDTH'd3846958;
publickey_row[5247] = `CIPHERTEXT_WIDTH'd11664961;
publickey_row[5248] = `CIPHERTEXT_WIDTH'd3914461;
publickey_row[5249] = `CIPHERTEXT_WIDTH'd4522773;
publickey_row[5250] = `CIPHERTEXT_WIDTH'd455533;
publickey_row[5251] = `CIPHERTEXT_WIDTH'd12303813;
publickey_row[5252] = `CIPHERTEXT_WIDTH'd3725991;
publickey_row[5253] = `CIPHERTEXT_WIDTH'd15201226;
publickey_row[5254] = `CIPHERTEXT_WIDTH'd12646074;
publickey_row[5255] = `CIPHERTEXT_WIDTH'd191387;
publickey_row[5256] = `CIPHERTEXT_WIDTH'd2769006;
publickey_row[5257] = `CIPHERTEXT_WIDTH'd3397000;
publickey_row[5258] = `CIPHERTEXT_WIDTH'd4920074;
publickey_row[5259] = `CIPHERTEXT_WIDTH'd5898261;
publickey_row[5260] = `CIPHERTEXT_WIDTH'd15726810;
publickey_row[5261] = `CIPHERTEXT_WIDTH'd9329568;
publickey_row[5262] = `CIPHERTEXT_WIDTH'd899470;
publickey_row[5263] = `CIPHERTEXT_WIDTH'd8241934;
publickey_row[5264] = `CIPHERTEXT_WIDTH'd7929330;
publickey_row[5265] = `CIPHERTEXT_WIDTH'd4180951;
publickey_row[5266] = `CIPHERTEXT_WIDTH'd8001035;
publickey_row[5267] = `CIPHERTEXT_WIDTH'd4377207;
publickey_row[5268] = `CIPHERTEXT_WIDTH'd12809945;
publickey_row[5269] = `CIPHERTEXT_WIDTH'd12104765;
publickey_row[5270] = `CIPHERTEXT_WIDTH'd11335807;
publickey_row[5271] = `CIPHERTEXT_WIDTH'd1937557;
publickey_row[5272] = `CIPHERTEXT_WIDTH'd6666453;
publickey_row[5273] = `CIPHERTEXT_WIDTH'd10550789;
publickey_row[5274] = `CIPHERTEXT_WIDTH'd1973007;
publickey_row[5275] = `CIPHERTEXT_WIDTH'd15137376;
publickey_row[5276] = `CIPHERTEXT_WIDTH'd5311632;
publickey_row[5277] = `CIPHERTEXT_WIDTH'd15857157;
publickey_row[5278] = `CIPHERTEXT_WIDTH'd13275428;
publickey_row[5279] = `CIPHERTEXT_WIDTH'd10890213;
publickey_row[5280] = `CIPHERTEXT_WIDTH'd11194262;
publickey_row[5281] = `CIPHERTEXT_WIDTH'd15765821;
publickey_row[5282] = `CIPHERTEXT_WIDTH'd9919155;
publickey_row[5283] = `CIPHERTEXT_WIDTH'd6526028;
publickey_row[5284] = `CIPHERTEXT_WIDTH'd11848454;
publickey_row[5285] = `CIPHERTEXT_WIDTH'd9562909;
publickey_row[5286] = `CIPHERTEXT_WIDTH'd3386336;
publickey_row[5287] = `CIPHERTEXT_WIDTH'd2974061;
publickey_row[5288] = `CIPHERTEXT_WIDTH'd7511540;
publickey_row[5289] = `CIPHERTEXT_WIDTH'd15265163;
publickey_row[5290] = `CIPHERTEXT_WIDTH'd9889696;
publickey_row[5291] = `CIPHERTEXT_WIDTH'd9956858;
publickey_row[5292] = `CIPHERTEXT_WIDTH'd2068390;
publickey_row[5293] = `CIPHERTEXT_WIDTH'd14591275;
publickey_row[5294] = `CIPHERTEXT_WIDTH'd6916570;
publickey_row[5295] = `CIPHERTEXT_WIDTH'd12540468;
publickey_row[5296] = `CIPHERTEXT_WIDTH'd13235147;
publickey_row[5297] = `CIPHERTEXT_WIDTH'd3996763;
publickey_row[5298] = `CIPHERTEXT_WIDTH'd11413824;
publickey_row[5299] = `CIPHERTEXT_WIDTH'd2474996;
publickey_row[5300] = `CIPHERTEXT_WIDTH'd7188407;
publickey_row[5301] = `CIPHERTEXT_WIDTH'd535553;
publickey_row[5302] = `CIPHERTEXT_WIDTH'd10916886;
publickey_row[5303] = `CIPHERTEXT_WIDTH'd11756609;
publickey_row[5304] = `CIPHERTEXT_WIDTH'd10102601;
publickey_row[5305] = `CIPHERTEXT_WIDTH'd15699867;
publickey_row[5306] = `CIPHERTEXT_WIDTH'd7044848;
publickey_row[5307] = `CIPHERTEXT_WIDTH'd6351237;
publickey_row[5308] = `CIPHERTEXT_WIDTH'd13322014;
publickey_row[5309] = `CIPHERTEXT_WIDTH'd3530368;
publickey_row[5310] = `CIPHERTEXT_WIDTH'd13005428;
publickey_row[5311] = `CIPHERTEXT_WIDTH'd5548053;
publickey_row[5312] = `CIPHERTEXT_WIDTH'd8641201;
publickey_row[5313] = `CIPHERTEXT_WIDTH'd11311342;
publickey_row[5314] = `CIPHERTEXT_WIDTH'd4593947;
publickey_row[5315] = `CIPHERTEXT_WIDTH'd16442148;
publickey_row[5316] = `CIPHERTEXT_WIDTH'd9311048;
publickey_row[5317] = `CIPHERTEXT_WIDTH'd726274;
publickey_row[5318] = `CIPHERTEXT_WIDTH'd16572538;
publickey_row[5319] = `CIPHERTEXT_WIDTH'd10656347;
publickey_row[5320] = `CIPHERTEXT_WIDTH'd345797;
publickey_row[5321] = `CIPHERTEXT_WIDTH'd4543352;
publickey_row[5322] = `CIPHERTEXT_WIDTH'd7165523;
publickey_row[5323] = `CIPHERTEXT_WIDTH'd230069;
publickey_row[5324] = `CIPHERTEXT_WIDTH'd10593820;
publickey_row[5325] = `CIPHERTEXT_WIDTH'd6447290;
publickey_row[5326] = `CIPHERTEXT_WIDTH'd3731786;
publickey_row[5327] = `CIPHERTEXT_WIDTH'd10718455;
publickey_row[5328] = `CIPHERTEXT_WIDTH'd9753953;
publickey_row[5329] = `CIPHERTEXT_WIDTH'd16472080;
publickey_row[5330] = `CIPHERTEXT_WIDTH'd10763822;
publickey_row[5331] = `CIPHERTEXT_WIDTH'd1161101;
publickey_row[5332] = `CIPHERTEXT_WIDTH'd12381651;
publickey_row[5333] = `CIPHERTEXT_WIDTH'd675739;
publickey_row[5334] = `CIPHERTEXT_WIDTH'd9401770;
publickey_row[5335] = `CIPHERTEXT_WIDTH'd66964;
publickey_row[5336] = `CIPHERTEXT_WIDTH'd4921294;
publickey_row[5337] = `CIPHERTEXT_WIDTH'd2185876;
publickey_row[5338] = `CIPHERTEXT_WIDTH'd4324394;
publickey_row[5339] = `CIPHERTEXT_WIDTH'd2834587;
publickey_row[5340] = `CIPHERTEXT_WIDTH'd6672493;
publickey_row[5341] = `CIPHERTEXT_WIDTH'd9136355;
publickey_row[5342] = `CIPHERTEXT_WIDTH'd15616692;
publickey_row[5343] = `CIPHERTEXT_WIDTH'd9865030;
publickey_row[5344] = `CIPHERTEXT_WIDTH'd5485780;
publickey_row[5345] = `CIPHERTEXT_WIDTH'd5438266;
publickey_row[5346] = `CIPHERTEXT_WIDTH'd6943126;
publickey_row[5347] = `CIPHERTEXT_WIDTH'd14060076;
publickey_row[5348] = `CIPHERTEXT_WIDTH'd12781941;
publickey_row[5349] = `CIPHERTEXT_WIDTH'd16380545;
publickey_row[5350] = `CIPHERTEXT_WIDTH'd6491557;
publickey_row[5351] = `CIPHERTEXT_WIDTH'd11939318;
publickey_row[5352] = `CIPHERTEXT_WIDTH'd15401543;
publickey_row[5353] = `CIPHERTEXT_WIDTH'd3121912;
publickey_row[5354] = `CIPHERTEXT_WIDTH'd15512514;
publickey_row[5355] = `CIPHERTEXT_WIDTH'd15504900;
publickey_row[5356] = `CIPHERTEXT_WIDTH'd14171144;
publickey_row[5357] = `CIPHERTEXT_WIDTH'd4314899;
publickey_row[5358] = `CIPHERTEXT_WIDTH'd14129592;
publickey_row[5359] = `CIPHERTEXT_WIDTH'd3106232;
publickey_row[5360] = `CIPHERTEXT_WIDTH'd11337833;
publickey_row[5361] = `CIPHERTEXT_WIDTH'd12643476;
publickey_row[5362] = `CIPHERTEXT_WIDTH'd10422173;
publickey_row[5363] = `CIPHERTEXT_WIDTH'd14231054;
publickey_row[5364] = `CIPHERTEXT_WIDTH'd2080369;
publickey_row[5365] = `CIPHERTEXT_WIDTH'd13505913;
publickey_row[5366] = `CIPHERTEXT_WIDTH'd4219240;
publickey_row[5367] = `CIPHERTEXT_WIDTH'd12318562;
publickey_row[5368] = `CIPHERTEXT_WIDTH'd2105485;
publickey_row[5369] = `CIPHERTEXT_WIDTH'd7294215;
publickey_row[5370] = `CIPHERTEXT_WIDTH'd3645510;
publickey_row[5371] = `CIPHERTEXT_WIDTH'd6961015;
publickey_row[5372] = `CIPHERTEXT_WIDTH'd1146014;
publickey_row[5373] = `CIPHERTEXT_WIDTH'd3170165;
publickey_row[5374] = `CIPHERTEXT_WIDTH'd4284074;
publickey_row[5375] = `CIPHERTEXT_WIDTH'd6273890;
publickey_row[5376] = `CIPHERTEXT_WIDTH'd11613216;
publickey_row[5377] = `CIPHERTEXT_WIDTH'd7530807;
publickey_row[5378] = `CIPHERTEXT_WIDTH'd9932348;
publickey_row[5379] = `CIPHERTEXT_WIDTH'd15851132;
publickey_row[5380] = `CIPHERTEXT_WIDTH'd2338895;
publickey_row[5381] = `CIPHERTEXT_WIDTH'd3419644;
publickey_row[5382] = `CIPHERTEXT_WIDTH'd10810016;
publickey_row[5383] = `CIPHERTEXT_WIDTH'd14682478;
publickey_row[5384] = `CIPHERTEXT_WIDTH'd5894613;
publickey_row[5385] = `CIPHERTEXT_WIDTH'd9244928;
publickey_row[5386] = `CIPHERTEXT_WIDTH'd15974583;
publickey_row[5387] = `CIPHERTEXT_WIDTH'd1249169;
publickey_row[5388] = `CIPHERTEXT_WIDTH'd9708049;
publickey_row[5389] = `CIPHERTEXT_WIDTH'd1544750;
publickey_row[5390] = `CIPHERTEXT_WIDTH'd4435263;
publickey_row[5391] = `CIPHERTEXT_WIDTH'd14065421;
publickey_row[5392] = `CIPHERTEXT_WIDTH'd2687586;
publickey_row[5393] = `CIPHERTEXT_WIDTH'd9686148;
publickey_row[5394] = `CIPHERTEXT_WIDTH'd4511306;
publickey_row[5395] = `CIPHERTEXT_WIDTH'd3653671;
publickey_row[5396] = `CIPHERTEXT_WIDTH'd15995538;
publickey_row[5397] = `CIPHERTEXT_WIDTH'd6201802;
publickey_row[5398] = `CIPHERTEXT_WIDTH'd6473888;
publickey_row[5399] = `CIPHERTEXT_WIDTH'd11535077;
publickey_row[5400] = `CIPHERTEXT_WIDTH'd1061657;
publickey_row[5401] = `CIPHERTEXT_WIDTH'd11166823;
publickey_row[5402] = `CIPHERTEXT_WIDTH'd14760151;
publickey_row[5403] = `CIPHERTEXT_WIDTH'd4789408;
publickey_row[5404] = `CIPHERTEXT_WIDTH'd2084420;
publickey_row[5405] = `CIPHERTEXT_WIDTH'd11098230;
publickey_row[5406] = `CIPHERTEXT_WIDTH'd1391220;
publickey_row[5407] = `CIPHERTEXT_WIDTH'd3822303;
publickey_row[5408] = `CIPHERTEXT_WIDTH'd9931314;
publickey_row[5409] = `CIPHERTEXT_WIDTH'd3783521;
publickey_row[5410] = `CIPHERTEXT_WIDTH'd324484;
publickey_row[5411] = `CIPHERTEXT_WIDTH'd8601229;
publickey_row[5412] = `CIPHERTEXT_WIDTH'd8836306;
publickey_row[5413] = `CIPHERTEXT_WIDTH'd1934845;
publickey_row[5414] = `CIPHERTEXT_WIDTH'd6677253;
publickey_row[5415] = `CIPHERTEXT_WIDTH'd5919391;
publickey_row[5416] = `CIPHERTEXT_WIDTH'd1028556;
publickey_row[5417] = `CIPHERTEXT_WIDTH'd1535028;
publickey_row[5418] = `CIPHERTEXT_WIDTH'd14484308;
publickey_row[5419] = `CIPHERTEXT_WIDTH'd5498489;
publickey_row[5420] = `CIPHERTEXT_WIDTH'd3622972;
publickey_row[5421] = `CIPHERTEXT_WIDTH'd15436690;
publickey_row[5422] = `CIPHERTEXT_WIDTH'd11902305;
publickey_row[5423] = `CIPHERTEXT_WIDTH'd11767046;
publickey_row[5424] = `CIPHERTEXT_WIDTH'd1616698;
publickey_row[5425] = `CIPHERTEXT_WIDTH'd253921;
publickey_row[5426] = `CIPHERTEXT_WIDTH'd10811037;
publickey_row[5427] = `CIPHERTEXT_WIDTH'd14884684;
publickey_row[5428] = `CIPHERTEXT_WIDTH'd364672;
publickey_row[5429] = `CIPHERTEXT_WIDTH'd11445370;
publickey_row[5430] = `CIPHERTEXT_WIDTH'd2013635;
publickey_row[5431] = `CIPHERTEXT_WIDTH'd919833;
publickey_row[5432] = `CIPHERTEXT_WIDTH'd9790871;
publickey_row[5433] = `CIPHERTEXT_WIDTH'd3972326;
publickey_row[5434] = `CIPHERTEXT_WIDTH'd3318990;
publickey_row[5435] = `CIPHERTEXT_WIDTH'd12132258;
publickey_row[5436] = `CIPHERTEXT_WIDTH'd9413565;
publickey_row[5437] = `CIPHERTEXT_WIDTH'd8468114;
publickey_row[5438] = `CIPHERTEXT_WIDTH'd13625438;
publickey_row[5439] = `CIPHERTEXT_WIDTH'd643809;
publickey_row[5440] = `CIPHERTEXT_WIDTH'd9643774;
publickey_row[5441] = `CIPHERTEXT_WIDTH'd11045491;
publickey_row[5442] = `CIPHERTEXT_WIDTH'd15171154;
publickey_row[5443] = `CIPHERTEXT_WIDTH'd15757452;
publickey_row[5444] = `CIPHERTEXT_WIDTH'd2495891;
publickey_row[5445] = `CIPHERTEXT_WIDTH'd2649222;
publickey_row[5446] = `CIPHERTEXT_WIDTH'd9495759;
publickey_row[5447] = `CIPHERTEXT_WIDTH'd3474734;
publickey_row[5448] = `CIPHERTEXT_WIDTH'd16585732;
publickey_row[5449] = `CIPHERTEXT_WIDTH'd10096019;
publickey_row[5450] = `CIPHERTEXT_WIDTH'd1847866;
publickey_row[5451] = `CIPHERTEXT_WIDTH'd7108901;
publickey_row[5452] = `CIPHERTEXT_WIDTH'd10926362;
publickey_row[5453] = `CIPHERTEXT_WIDTH'd890706;
publickey_row[5454] = `CIPHERTEXT_WIDTH'd1027554;
publickey_row[5455] = `CIPHERTEXT_WIDTH'd12010500;
publickey_row[5456] = `CIPHERTEXT_WIDTH'd3665956;
publickey_row[5457] = `CIPHERTEXT_WIDTH'd774302;
publickey_row[5458] = `CIPHERTEXT_WIDTH'd10893024;
publickey_row[5459] = `CIPHERTEXT_WIDTH'd9673997;
publickey_row[5460] = `CIPHERTEXT_WIDTH'd1579153;
publickey_row[5461] = `CIPHERTEXT_WIDTH'd1800761;
publickey_row[5462] = `CIPHERTEXT_WIDTH'd12062582;
publickey_row[5463] = `CIPHERTEXT_WIDTH'd15300956;
publickey_row[5464] = `CIPHERTEXT_WIDTH'd16241243;
publickey_row[5465] = `CIPHERTEXT_WIDTH'd2890251;
publickey_row[5466] = `CIPHERTEXT_WIDTH'd3637139;
publickey_row[5467] = `CIPHERTEXT_WIDTH'd14984680;
publickey_row[5468] = `CIPHERTEXT_WIDTH'd5691365;
publickey_row[5469] = `CIPHERTEXT_WIDTH'd296536;
publickey_row[5470] = `CIPHERTEXT_WIDTH'd13719106;
publickey_row[5471] = `CIPHERTEXT_WIDTH'd7679491;
publickey_row[5472] = `CIPHERTEXT_WIDTH'd12144061;
publickey_row[5473] = `CIPHERTEXT_WIDTH'd1595429;
publickey_row[5474] = `CIPHERTEXT_WIDTH'd10231954;
publickey_row[5475] = `CIPHERTEXT_WIDTH'd5950291;
publickey_row[5476] = `CIPHERTEXT_WIDTH'd7514001;
publickey_row[5477] = `CIPHERTEXT_WIDTH'd4714256;
publickey_row[5478] = `CIPHERTEXT_WIDTH'd14663799;
publickey_row[5479] = `CIPHERTEXT_WIDTH'd16460278;
publickey_row[5480] = `CIPHERTEXT_WIDTH'd13936377;
publickey_row[5481] = `CIPHERTEXT_WIDTH'd6486007;
publickey_row[5482] = `CIPHERTEXT_WIDTH'd11828826;
publickey_row[5483] = `CIPHERTEXT_WIDTH'd10331141;
publickey_row[5484] = `CIPHERTEXT_WIDTH'd12644952;
publickey_row[5485] = `CIPHERTEXT_WIDTH'd8195679;
publickey_row[5486] = `CIPHERTEXT_WIDTH'd998344;
publickey_row[5487] = `CIPHERTEXT_WIDTH'd6643637;
publickey_row[5488] = `CIPHERTEXT_WIDTH'd13005460;
publickey_row[5489] = `CIPHERTEXT_WIDTH'd13852355;
publickey_row[5490] = `CIPHERTEXT_WIDTH'd11147912;
publickey_row[5491] = `CIPHERTEXT_WIDTH'd3609018;
publickey_row[5492] = `CIPHERTEXT_WIDTH'd5614394;
publickey_row[5493] = `CIPHERTEXT_WIDTH'd13111289;
publickey_row[5494] = `CIPHERTEXT_WIDTH'd6771989;
publickey_row[5495] = `CIPHERTEXT_WIDTH'd8924716;
publickey_row[5496] = `CIPHERTEXT_WIDTH'd12871918;
publickey_row[5497] = `CIPHERTEXT_WIDTH'd4185374;
publickey_row[5498] = `CIPHERTEXT_WIDTH'd346648;
publickey_row[5499] = `CIPHERTEXT_WIDTH'd5896949;
publickey_row[5500] = `CIPHERTEXT_WIDTH'd10605031;
publickey_row[5501] = `CIPHERTEXT_WIDTH'd8820483;
publickey_row[5502] = `CIPHERTEXT_WIDTH'd3797997;
publickey_row[5503] = `CIPHERTEXT_WIDTH'd9878478;
publickey_row[5504] = `CIPHERTEXT_WIDTH'd12607263;
publickey_row[5505] = `CIPHERTEXT_WIDTH'd14711252;
publickey_row[5506] = `CIPHERTEXT_WIDTH'd7268505;
publickey_row[5507] = `CIPHERTEXT_WIDTH'd7241141;
publickey_row[5508] = `CIPHERTEXT_WIDTH'd14347180;
publickey_row[5509] = `CIPHERTEXT_WIDTH'd16047596;
publickey_row[5510] = `CIPHERTEXT_WIDTH'd8784227;
publickey_row[5511] = `CIPHERTEXT_WIDTH'd5916187;
publickey_row[5512] = `CIPHERTEXT_WIDTH'd6770709;
publickey_row[5513] = `CIPHERTEXT_WIDTH'd7087477;
publickey_row[5514] = `CIPHERTEXT_WIDTH'd3335254;
publickey_row[5515] = `CIPHERTEXT_WIDTH'd4010810;
publickey_row[5516] = `CIPHERTEXT_WIDTH'd9152265;
publickey_row[5517] = `CIPHERTEXT_WIDTH'd16117485;
publickey_row[5518] = `CIPHERTEXT_WIDTH'd6020700;
publickey_row[5519] = `CIPHERTEXT_WIDTH'd12833887;
publickey_row[5520] = `CIPHERTEXT_WIDTH'd7940064;
publickey_row[5521] = `CIPHERTEXT_WIDTH'd9273786;
publickey_row[5522] = `CIPHERTEXT_WIDTH'd9998380;
publickey_row[5523] = `CIPHERTEXT_WIDTH'd5523278;
publickey_row[5524] = `CIPHERTEXT_WIDTH'd6456210;
publickey_row[5525] = `CIPHERTEXT_WIDTH'd14781771;
publickey_row[5526] = `CIPHERTEXT_WIDTH'd6464436;
publickey_row[5527] = `CIPHERTEXT_WIDTH'd9228546;
publickey_row[5528] = `CIPHERTEXT_WIDTH'd10206839;
publickey_row[5529] = `CIPHERTEXT_WIDTH'd8703228;
publickey_row[5530] = `CIPHERTEXT_WIDTH'd7114556;
publickey_row[5531] = `CIPHERTEXT_WIDTH'd4736791;
publickey_row[5532] = `CIPHERTEXT_WIDTH'd15964460;
publickey_row[5533] = `CIPHERTEXT_WIDTH'd1614012;
publickey_row[5534] = `CIPHERTEXT_WIDTH'd7040851;
publickey_row[5535] = `CIPHERTEXT_WIDTH'd14870732;
publickey_row[5536] = `CIPHERTEXT_WIDTH'd9561002;
publickey_row[5537] = `CIPHERTEXT_WIDTH'd8569725;
publickey_row[5538] = `CIPHERTEXT_WIDTH'd6217738;
publickey_row[5539] = `CIPHERTEXT_WIDTH'd12433923;
publickey_row[5540] = `CIPHERTEXT_WIDTH'd4325062;
publickey_row[5541] = `CIPHERTEXT_WIDTH'd6934048;
publickey_row[5542] = `CIPHERTEXT_WIDTH'd14347724;
publickey_row[5543] = `CIPHERTEXT_WIDTH'd6940654;
publickey_row[5544] = `CIPHERTEXT_WIDTH'd15081254;
publickey_row[5545] = `CIPHERTEXT_WIDTH'd16497339;
publickey_row[5546] = `CIPHERTEXT_WIDTH'd14508833;
publickey_row[5547] = `CIPHERTEXT_WIDTH'd12012657;
publickey_row[5548] = `CIPHERTEXT_WIDTH'd14076003;
publickey_row[5549] = `CIPHERTEXT_WIDTH'd9558006;
publickey_row[5550] = `CIPHERTEXT_WIDTH'd279803;
publickey_row[5551] = `CIPHERTEXT_WIDTH'd5312088;
publickey_row[5552] = `CIPHERTEXT_WIDTH'd5927626;
publickey_row[5553] = `CIPHERTEXT_WIDTH'd3785438;
publickey_row[5554] = `CIPHERTEXT_WIDTH'd7129967;
publickey_row[5555] = `CIPHERTEXT_WIDTH'd16611282;
publickey_row[5556] = `CIPHERTEXT_WIDTH'd9935323;
publickey_row[5557] = `CIPHERTEXT_WIDTH'd8450529;
publickey_row[5558] = `CIPHERTEXT_WIDTH'd10937112;
publickey_row[5559] = `CIPHERTEXT_WIDTH'd10807623;
publickey_row[5560] = `CIPHERTEXT_WIDTH'd5452036;
publickey_row[5561] = `CIPHERTEXT_WIDTH'd13450038;
publickey_row[5562] = `CIPHERTEXT_WIDTH'd13294872;
publickey_row[5563] = `CIPHERTEXT_WIDTH'd6424387;
publickey_row[5564] = `CIPHERTEXT_WIDTH'd16466640;
publickey_row[5565] = `CIPHERTEXT_WIDTH'd15910262;
publickey_row[5566] = `CIPHERTEXT_WIDTH'd5414665;
publickey_row[5567] = `CIPHERTEXT_WIDTH'd3025748;
publickey_row[5568] = `CIPHERTEXT_WIDTH'd9604834;
publickey_row[5569] = `CIPHERTEXT_WIDTH'd11740913;
publickey_row[5570] = `CIPHERTEXT_WIDTH'd1029128;
publickey_row[5571] = `CIPHERTEXT_WIDTH'd13195353;
publickey_row[5572] = `CIPHERTEXT_WIDTH'd16740272;
publickey_row[5573] = `CIPHERTEXT_WIDTH'd11530922;
publickey_row[5574] = `CIPHERTEXT_WIDTH'd3399634;
publickey_row[5575] = `CIPHERTEXT_WIDTH'd4070103;
publickey_row[5576] = `CIPHERTEXT_WIDTH'd7994509;
publickey_row[5577] = `CIPHERTEXT_WIDTH'd11702334;
publickey_row[5578] = `CIPHERTEXT_WIDTH'd10079337;
publickey_row[5579] = `CIPHERTEXT_WIDTH'd11745532;
publickey_row[5580] = `CIPHERTEXT_WIDTH'd14909664;
publickey_row[5581] = `CIPHERTEXT_WIDTH'd12174832;
publickey_row[5582] = `CIPHERTEXT_WIDTH'd6356234;
publickey_row[5583] = `CIPHERTEXT_WIDTH'd13815480;
publickey_row[5584] = `CIPHERTEXT_WIDTH'd12659988;
publickey_row[5585] = `CIPHERTEXT_WIDTH'd15045340;
publickey_row[5586] = `CIPHERTEXT_WIDTH'd13486105;
publickey_row[5587] = `CIPHERTEXT_WIDTH'd1049417;
publickey_row[5588] = `CIPHERTEXT_WIDTH'd1014485;
publickey_row[5589] = `CIPHERTEXT_WIDTH'd6293540;
publickey_row[5590] = `CIPHERTEXT_WIDTH'd3989932;
publickey_row[5591] = `CIPHERTEXT_WIDTH'd12538493;
publickey_row[5592] = `CIPHERTEXT_WIDTH'd11295568;
publickey_row[5593] = `CIPHERTEXT_WIDTH'd16505307;
publickey_row[5594] = `CIPHERTEXT_WIDTH'd16702502;
publickey_row[5595] = `CIPHERTEXT_WIDTH'd5283439;
publickey_row[5596] = `CIPHERTEXT_WIDTH'd483252;
publickey_row[5597] = `CIPHERTEXT_WIDTH'd8249333;
publickey_row[5598] = `CIPHERTEXT_WIDTH'd8775888;
publickey_row[5599] = `CIPHERTEXT_WIDTH'd14390823;
publickey_row[5600] = `CIPHERTEXT_WIDTH'd7908285;
publickey_row[5601] = `CIPHERTEXT_WIDTH'd13142267;
publickey_row[5602] = `CIPHERTEXT_WIDTH'd11722272;
publickey_row[5603] = `CIPHERTEXT_WIDTH'd14608003;
publickey_row[5604] = `CIPHERTEXT_WIDTH'd14341404;
publickey_row[5605] = `CIPHERTEXT_WIDTH'd2653258;
publickey_row[5606] = `CIPHERTEXT_WIDTH'd13012363;
publickey_row[5607] = `CIPHERTEXT_WIDTH'd5414035;
publickey_row[5608] = `CIPHERTEXT_WIDTH'd13122067;
publickey_row[5609] = `CIPHERTEXT_WIDTH'd2806997;
publickey_row[5610] = `CIPHERTEXT_WIDTH'd12719692;
publickey_row[5611] = `CIPHERTEXT_WIDTH'd8222084;
publickey_row[5612] = `CIPHERTEXT_WIDTH'd14539958;
publickey_row[5613] = `CIPHERTEXT_WIDTH'd16337097;
publickey_row[5614] = `CIPHERTEXT_WIDTH'd9709181;
publickey_row[5615] = `CIPHERTEXT_WIDTH'd749199;
publickey_row[5616] = `CIPHERTEXT_WIDTH'd9055996;
publickey_row[5617] = `CIPHERTEXT_WIDTH'd13670384;
publickey_row[5618] = `CIPHERTEXT_WIDTH'd13361751;
publickey_row[5619] = `CIPHERTEXT_WIDTH'd3264356;
publickey_row[5620] = `CIPHERTEXT_WIDTH'd15279453;
publickey_row[5621] = `CIPHERTEXT_WIDTH'd6280520;
publickey_row[5622] = `CIPHERTEXT_WIDTH'd16037529;
publickey_row[5623] = `CIPHERTEXT_WIDTH'd15975477;
publickey_row[5624] = `CIPHERTEXT_WIDTH'd13124666;
publickey_row[5625] = `CIPHERTEXT_WIDTH'd1492972;
publickey_row[5626] = `CIPHERTEXT_WIDTH'd1066370;
publickey_row[5627] = `CIPHERTEXT_WIDTH'd7975718;
publickey_row[5628] = `CIPHERTEXT_WIDTH'd766276;
publickey_row[5629] = `CIPHERTEXT_WIDTH'd10532117;
publickey_row[5630] = `CIPHERTEXT_WIDTH'd4162265;
publickey_row[5631] = `CIPHERTEXT_WIDTH'd5773436;
publickey_row[5632] = `CIPHERTEXT_WIDTH'd2234062;
publickey_row[5633] = `CIPHERTEXT_WIDTH'd8311537;
publickey_row[5634] = `CIPHERTEXT_WIDTH'd11844788;
publickey_row[5635] = `CIPHERTEXT_WIDTH'd10215943;
publickey_row[5636] = `CIPHERTEXT_WIDTH'd12546528;
publickey_row[5637] = `CIPHERTEXT_WIDTH'd9535304;
publickey_row[5638] = `CIPHERTEXT_WIDTH'd124662;
publickey_row[5639] = `CIPHERTEXT_WIDTH'd12559585;
publickey_row[5640] = `CIPHERTEXT_WIDTH'd14142061;
publickey_row[5641] = `CIPHERTEXT_WIDTH'd10011540;
publickey_row[5642] = `CIPHERTEXT_WIDTH'd4644395;
publickey_row[5643] = `CIPHERTEXT_WIDTH'd14163073;
publickey_row[5644] = `CIPHERTEXT_WIDTH'd4835231;
publickey_row[5645] = `CIPHERTEXT_WIDTH'd16152019;
publickey_row[5646] = `CIPHERTEXT_WIDTH'd8806850;
publickey_row[5647] = `CIPHERTEXT_WIDTH'd6315257;
publickey_row[5648] = `CIPHERTEXT_WIDTH'd7370835;
publickey_row[5649] = `CIPHERTEXT_WIDTH'd7284106;
publickey_row[5650] = `CIPHERTEXT_WIDTH'd7194570;
publickey_row[5651] = `CIPHERTEXT_WIDTH'd699715;
publickey_row[5652] = `CIPHERTEXT_WIDTH'd58758;
publickey_row[5653] = `CIPHERTEXT_WIDTH'd152826;
publickey_row[5654] = `CIPHERTEXT_WIDTH'd7412769;
publickey_row[5655] = `CIPHERTEXT_WIDTH'd13185330;
publickey_row[5656] = `CIPHERTEXT_WIDTH'd3310265;
publickey_row[5657] = `CIPHERTEXT_WIDTH'd7393683;
publickey_row[5658] = `CIPHERTEXT_WIDTH'd13069352;
publickey_row[5659] = `CIPHERTEXT_WIDTH'd13562324;
publickey_row[5660] = `CIPHERTEXT_WIDTH'd10393996;
publickey_row[5661] = `CIPHERTEXT_WIDTH'd7647303;
publickey_row[5662] = `CIPHERTEXT_WIDTH'd12081858;
publickey_row[5663] = `CIPHERTEXT_WIDTH'd15727558;
publickey_row[5664] = `CIPHERTEXT_WIDTH'd4737441;
publickey_row[5665] = `CIPHERTEXT_WIDTH'd1055593;
publickey_row[5666] = `CIPHERTEXT_WIDTH'd6423904;
publickey_row[5667] = `CIPHERTEXT_WIDTH'd1595199;
publickey_row[5668] = `CIPHERTEXT_WIDTH'd13115548;
publickey_row[5669] = `CIPHERTEXT_WIDTH'd6928797;
publickey_row[5670] = `CIPHERTEXT_WIDTH'd5701385;
publickey_row[5671] = `CIPHERTEXT_WIDTH'd10222283;
publickey_row[5672] = `CIPHERTEXT_WIDTH'd3974871;
publickey_row[5673] = `CIPHERTEXT_WIDTH'd10409787;
publickey_row[5674] = `CIPHERTEXT_WIDTH'd13782350;
publickey_row[5675] = `CIPHERTEXT_WIDTH'd15776762;
publickey_row[5676] = `CIPHERTEXT_WIDTH'd12153450;
publickey_row[5677] = `CIPHERTEXT_WIDTH'd13980075;
publickey_row[5678] = `CIPHERTEXT_WIDTH'd198767;
publickey_row[5679] = `CIPHERTEXT_WIDTH'd664782;
publickey_row[5680] = `CIPHERTEXT_WIDTH'd3051289;
publickey_row[5681] = `CIPHERTEXT_WIDTH'd15435574;
publickey_row[5682] = `CIPHERTEXT_WIDTH'd3440671;
publickey_row[5683] = `CIPHERTEXT_WIDTH'd15218865;
publickey_row[5684] = `CIPHERTEXT_WIDTH'd2068954;
publickey_row[5685] = `CIPHERTEXT_WIDTH'd8834375;
publickey_row[5686] = `CIPHERTEXT_WIDTH'd4407165;
publickey_row[5687] = `CIPHERTEXT_WIDTH'd5004656;
publickey_row[5688] = `CIPHERTEXT_WIDTH'd5938971;
publickey_row[5689] = `CIPHERTEXT_WIDTH'd3011659;
publickey_row[5690] = `CIPHERTEXT_WIDTH'd12153091;
publickey_row[5691] = `CIPHERTEXT_WIDTH'd14564547;
publickey_row[5692] = `CIPHERTEXT_WIDTH'd11431231;
publickey_row[5693] = `CIPHERTEXT_WIDTH'd2122593;
publickey_row[5694] = `CIPHERTEXT_WIDTH'd9724584;
publickey_row[5695] = `CIPHERTEXT_WIDTH'd11813965;
publickey_row[5696] = `CIPHERTEXT_WIDTH'd13981747;
publickey_row[5697] = `CIPHERTEXT_WIDTH'd7789691;
publickey_row[5698] = `CIPHERTEXT_WIDTH'd6642503;
publickey_row[5699] = `CIPHERTEXT_WIDTH'd4523180;
publickey_row[5700] = `CIPHERTEXT_WIDTH'd9425729;
publickey_row[5701] = `CIPHERTEXT_WIDTH'd3971129;
publickey_row[5702] = `CIPHERTEXT_WIDTH'd15882567;
publickey_row[5703] = `CIPHERTEXT_WIDTH'd5617055;
publickey_row[5704] = `CIPHERTEXT_WIDTH'd13248883;
publickey_row[5705] = `CIPHERTEXT_WIDTH'd1314641;
publickey_row[5706] = `CIPHERTEXT_WIDTH'd8496579;
publickey_row[5707] = `CIPHERTEXT_WIDTH'd10489865;
publickey_row[5708] = `CIPHERTEXT_WIDTH'd3705130;
publickey_row[5709] = `CIPHERTEXT_WIDTH'd1960065;
publickey_row[5710] = `CIPHERTEXT_WIDTH'd9832436;
publickey_row[5711] = `CIPHERTEXT_WIDTH'd13453336;
publickey_row[5712] = `CIPHERTEXT_WIDTH'd9850193;
publickey_row[5713] = `CIPHERTEXT_WIDTH'd350761;
publickey_row[5714] = `CIPHERTEXT_WIDTH'd3929308;
publickey_row[5715] = `CIPHERTEXT_WIDTH'd12843522;
publickey_row[5716] = `CIPHERTEXT_WIDTH'd9215507;
publickey_row[5717] = `CIPHERTEXT_WIDTH'd10668386;
publickey_row[5718] = `CIPHERTEXT_WIDTH'd4386214;
publickey_row[5719] = `CIPHERTEXT_WIDTH'd14568431;
publickey_row[5720] = `CIPHERTEXT_WIDTH'd1622010;
publickey_row[5721] = `CIPHERTEXT_WIDTH'd15827783;
publickey_row[5722] = `CIPHERTEXT_WIDTH'd6705887;
publickey_row[5723] = `CIPHERTEXT_WIDTH'd10737744;
publickey_row[5724] = `CIPHERTEXT_WIDTH'd1954041;
publickey_row[5725] = `CIPHERTEXT_WIDTH'd6463730;
publickey_row[5726] = `CIPHERTEXT_WIDTH'd2696275;
publickey_row[5727] = `CIPHERTEXT_WIDTH'd12857951;
publickey_row[5728] = `CIPHERTEXT_WIDTH'd3636830;
publickey_row[5729] = `CIPHERTEXT_WIDTH'd14972979;
publickey_row[5730] = `CIPHERTEXT_WIDTH'd15870358;
publickey_row[5731] = `CIPHERTEXT_WIDTH'd16553337;
publickey_row[5732] = `CIPHERTEXT_WIDTH'd15097953;
publickey_row[5733] = `CIPHERTEXT_WIDTH'd11751361;
publickey_row[5734] = `CIPHERTEXT_WIDTH'd2090234;
publickey_row[5735] = `CIPHERTEXT_WIDTH'd5322159;
publickey_row[5736] = `CIPHERTEXT_WIDTH'd12320084;
publickey_row[5737] = `CIPHERTEXT_WIDTH'd12821233;
publickey_row[5738] = `CIPHERTEXT_WIDTH'd12140666;
publickey_row[5739] = `CIPHERTEXT_WIDTH'd8367631;
publickey_row[5740] = `CIPHERTEXT_WIDTH'd7232133;
publickey_row[5741] = `CIPHERTEXT_WIDTH'd11925771;
publickey_row[5742] = `CIPHERTEXT_WIDTH'd790546;
publickey_row[5743] = `CIPHERTEXT_WIDTH'd16210215;
publickey_row[5744] = `CIPHERTEXT_WIDTH'd15693456;
publickey_row[5745] = `CIPHERTEXT_WIDTH'd11381416;
publickey_row[5746] = `CIPHERTEXT_WIDTH'd5830751;
publickey_row[5747] = `CIPHERTEXT_WIDTH'd7396597;
publickey_row[5748] = `CIPHERTEXT_WIDTH'd2862213;
publickey_row[5749] = `CIPHERTEXT_WIDTH'd13035642;
publickey_row[5750] = `CIPHERTEXT_WIDTH'd5517871;
publickey_row[5751] = `CIPHERTEXT_WIDTH'd3087317;
publickey_row[5752] = `CIPHERTEXT_WIDTH'd13909121;
publickey_row[5753] = `CIPHERTEXT_WIDTH'd10098308;
publickey_row[5754] = `CIPHERTEXT_WIDTH'd5561311;
publickey_row[5755] = `CIPHERTEXT_WIDTH'd1378843;
publickey_row[5756] = `CIPHERTEXT_WIDTH'd9526686;
publickey_row[5757] = `CIPHERTEXT_WIDTH'd6549408;
publickey_row[5758] = `CIPHERTEXT_WIDTH'd1023514;
publickey_row[5759] = `CIPHERTEXT_WIDTH'd14296718;
publickey_row[5760] = `CIPHERTEXT_WIDTH'd6254071;
publickey_row[5761] = `CIPHERTEXT_WIDTH'd8739990;
publickey_row[5762] = `CIPHERTEXT_WIDTH'd4657556;
publickey_row[5763] = `CIPHERTEXT_WIDTH'd9401207;
publickey_row[5764] = `CIPHERTEXT_WIDTH'd1750749;
publickey_row[5765] = `CIPHERTEXT_WIDTH'd5347612;
publickey_row[5766] = `CIPHERTEXT_WIDTH'd8324183;
publickey_row[5767] = `CIPHERTEXT_WIDTH'd5469038;
publickey_row[5768] = `CIPHERTEXT_WIDTH'd9348436;
publickey_row[5769] = `CIPHERTEXT_WIDTH'd5439300;
publickey_row[5770] = `CIPHERTEXT_WIDTH'd12611793;
publickey_row[5771] = `CIPHERTEXT_WIDTH'd4192964;
publickey_row[5772] = `CIPHERTEXT_WIDTH'd2682368;
publickey_row[5773] = `CIPHERTEXT_WIDTH'd13947129;
publickey_row[5774] = `CIPHERTEXT_WIDTH'd15481532;
publickey_row[5775] = `CIPHERTEXT_WIDTH'd15760178;
publickey_row[5776] = `CIPHERTEXT_WIDTH'd14777667;
publickey_row[5777] = `CIPHERTEXT_WIDTH'd9360061;
publickey_row[5778] = `CIPHERTEXT_WIDTH'd3437042;
publickey_row[5779] = `CIPHERTEXT_WIDTH'd8812814;
publickey_row[5780] = `CIPHERTEXT_WIDTH'd2972907;
publickey_row[5781] = `CIPHERTEXT_WIDTH'd11219189;
publickey_row[5782] = `CIPHERTEXT_WIDTH'd10267507;
publickey_row[5783] = `CIPHERTEXT_WIDTH'd624413;
publickey_row[5784] = `CIPHERTEXT_WIDTH'd5540272;
publickey_row[5785] = `CIPHERTEXT_WIDTH'd1823463;
publickey_row[5786] = `CIPHERTEXT_WIDTH'd11145042;
publickey_row[5787] = `CIPHERTEXT_WIDTH'd6906916;
publickey_row[5788] = `CIPHERTEXT_WIDTH'd5896510;
publickey_row[5789] = `CIPHERTEXT_WIDTH'd2359159;
publickey_row[5790] = `CIPHERTEXT_WIDTH'd6359185;
publickey_row[5791] = `CIPHERTEXT_WIDTH'd9250347;
publickey_row[5792] = `CIPHERTEXT_WIDTH'd11756594;
publickey_row[5793] = `CIPHERTEXT_WIDTH'd13825751;
publickey_row[5794] = `CIPHERTEXT_WIDTH'd4612912;
publickey_row[5795] = `CIPHERTEXT_WIDTH'd10743777;
publickey_row[5796] = `CIPHERTEXT_WIDTH'd1672065;
publickey_row[5797] = `CIPHERTEXT_WIDTH'd4272028;
publickey_row[5798] = `CIPHERTEXT_WIDTH'd7518803;
publickey_row[5799] = `CIPHERTEXT_WIDTH'd1722670;
publickey_row[5800] = `CIPHERTEXT_WIDTH'd6165161;
publickey_row[5801] = `CIPHERTEXT_WIDTH'd6333031;
publickey_row[5802] = `CIPHERTEXT_WIDTH'd2512372;
publickey_row[5803] = `CIPHERTEXT_WIDTH'd3844675;
publickey_row[5804] = `CIPHERTEXT_WIDTH'd5214031;
publickey_row[5805] = `CIPHERTEXT_WIDTH'd14795377;
publickey_row[5806] = `CIPHERTEXT_WIDTH'd3261329;
publickey_row[5807] = `CIPHERTEXT_WIDTH'd14285269;
publickey_row[5808] = `CIPHERTEXT_WIDTH'd7834118;
publickey_row[5809] = `CIPHERTEXT_WIDTH'd7734201;
publickey_row[5810] = `CIPHERTEXT_WIDTH'd3147302;
publickey_row[5811] = `CIPHERTEXT_WIDTH'd16682445;
publickey_row[5812] = `CIPHERTEXT_WIDTH'd7175110;
publickey_row[5813] = `CIPHERTEXT_WIDTH'd13568034;
publickey_row[5814] = `CIPHERTEXT_WIDTH'd14134260;
publickey_row[5815] = `CIPHERTEXT_WIDTH'd9655025;
publickey_row[5816] = `CIPHERTEXT_WIDTH'd2871567;
publickey_row[5817] = `CIPHERTEXT_WIDTH'd3338926;
publickey_row[5818] = `CIPHERTEXT_WIDTH'd12343987;
publickey_row[5819] = `CIPHERTEXT_WIDTH'd15929296;
publickey_row[5820] = `CIPHERTEXT_WIDTH'd13335705;
publickey_row[5821] = `CIPHERTEXT_WIDTH'd10035321;
publickey_row[5822] = `CIPHERTEXT_WIDTH'd8702741;
publickey_row[5823] = `CIPHERTEXT_WIDTH'd706313;
publickey_row[5824] = `CIPHERTEXT_WIDTH'd458664;
publickey_row[5825] = `CIPHERTEXT_WIDTH'd9785512;
publickey_row[5826] = `CIPHERTEXT_WIDTH'd3904762;
publickey_row[5827] = `CIPHERTEXT_WIDTH'd2760341;
publickey_row[5828] = `CIPHERTEXT_WIDTH'd5811119;
publickey_row[5829] = `CIPHERTEXT_WIDTH'd3246702;
publickey_row[5830] = `CIPHERTEXT_WIDTH'd16226450;
publickey_row[5831] = `CIPHERTEXT_WIDTH'd319933;
publickey_row[5832] = `CIPHERTEXT_WIDTH'd14817639;
publickey_row[5833] = `CIPHERTEXT_WIDTH'd14066615;
publickey_row[5834] = `CIPHERTEXT_WIDTH'd555967;
publickey_row[5835] = `CIPHERTEXT_WIDTH'd12435352;
publickey_row[5836] = `CIPHERTEXT_WIDTH'd7353788;
publickey_row[5837] = `CIPHERTEXT_WIDTH'd15158426;
publickey_row[5838] = `CIPHERTEXT_WIDTH'd12642787;
publickey_row[5839] = `CIPHERTEXT_WIDTH'd10025213;
publickey_row[5840] = `CIPHERTEXT_WIDTH'd2953435;
publickey_row[5841] = `CIPHERTEXT_WIDTH'd13622490;
publickey_row[5842] = `CIPHERTEXT_WIDTH'd10695175;
publickey_row[5843] = `CIPHERTEXT_WIDTH'd15081692;
publickey_row[5844] = `CIPHERTEXT_WIDTH'd16774;
publickey_row[5845] = `CIPHERTEXT_WIDTH'd6606887;
publickey_row[5846] = `CIPHERTEXT_WIDTH'd7989956;
publickey_row[5847] = `CIPHERTEXT_WIDTH'd9098601;
publickey_row[5848] = `CIPHERTEXT_WIDTH'd13568019;
publickey_row[5849] = `CIPHERTEXT_WIDTH'd3511577;
publickey_row[5850] = `CIPHERTEXT_WIDTH'd3643284;
publickey_row[5851] = `CIPHERTEXT_WIDTH'd534561;
publickey_row[5852] = `CIPHERTEXT_WIDTH'd9175522;
publickey_row[5853] = `CIPHERTEXT_WIDTH'd8856491;
publickey_row[5854] = `CIPHERTEXT_WIDTH'd1102895;
publickey_row[5855] = `CIPHERTEXT_WIDTH'd9711842;
publickey_row[5856] = `CIPHERTEXT_WIDTH'd13627419;
publickey_row[5857] = `CIPHERTEXT_WIDTH'd16407536;
publickey_row[5858] = `CIPHERTEXT_WIDTH'd803194;
publickey_row[5859] = `CIPHERTEXT_WIDTH'd11646597;
publickey_row[5860] = `CIPHERTEXT_WIDTH'd8709968;
publickey_row[5861] = `CIPHERTEXT_WIDTH'd8284557;
publickey_row[5862] = `CIPHERTEXT_WIDTH'd16057636;
publickey_row[5863] = `CIPHERTEXT_WIDTH'd5285491;
publickey_row[5864] = `CIPHERTEXT_WIDTH'd1258376;
publickey_row[5865] = `CIPHERTEXT_WIDTH'd4783259;
publickey_row[5866] = `CIPHERTEXT_WIDTH'd11979286;
publickey_row[5867] = `CIPHERTEXT_WIDTH'd13808379;
publickey_row[5868] = `CIPHERTEXT_WIDTH'd11282563;
publickey_row[5869] = `CIPHERTEXT_WIDTH'd13710543;
publickey_row[5870] = `CIPHERTEXT_WIDTH'd11142332;
publickey_row[5871] = `CIPHERTEXT_WIDTH'd15572291;
publickey_row[5872] = `CIPHERTEXT_WIDTH'd7506832;
publickey_row[5873] = `CIPHERTEXT_WIDTH'd2838939;
publickey_row[5874] = `CIPHERTEXT_WIDTH'd3275024;
publickey_row[5875] = `CIPHERTEXT_WIDTH'd11627291;
publickey_row[5876] = `CIPHERTEXT_WIDTH'd14104109;
publickey_row[5877] = `CIPHERTEXT_WIDTH'd3788890;
publickey_row[5878] = `CIPHERTEXT_WIDTH'd11820408;
publickey_row[5879] = `CIPHERTEXT_WIDTH'd7030037;
publickey_row[5880] = `CIPHERTEXT_WIDTH'd14298449;
publickey_row[5881] = `CIPHERTEXT_WIDTH'd608086;
publickey_row[5882] = `CIPHERTEXT_WIDTH'd3283847;
publickey_row[5883] = `CIPHERTEXT_WIDTH'd13347517;
publickey_row[5884] = `CIPHERTEXT_WIDTH'd12172463;
publickey_row[5885] = `CIPHERTEXT_WIDTH'd15065809;
publickey_row[5886] = `CIPHERTEXT_WIDTH'd12176056;
publickey_row[5887] = `CIPHERTEXT_WIDTH'd3154858;
publickey_row[5888] = `CIPHERTEXT_WIDTH'd4856128;
publickey_row[5889] = `CIPHERTEXT_WIDTH'd4827007;
publickey_row[5890] = `CIPHERTEXT_WIDTH'd4111247;
publickey_row[5891] = `CIPHERTEXT_WIDTH'd5516055;
publickey_row[5892] = `CIPHERTEXT_WIDTH'd5378527;
publickey_row[5893] = `CIPHERTEXT_WIDTH'd15463665;
publickey_row[5894] = `CIPHERTEXT_WIDTH'd14848460;
publickey_row[5895] = `CIPHERTEXT_WIDTH'd4984057;
publickey_row[5896] = `CIPHERTEXT_WIDTH'd4180784;
publickey_row[5897] = `CIPHERTEXT_WIDTH'd8388794;
publickey_row[5898] = `CIPHERTEXT_WIDTH'd5621040;
publickey_row[5899] = `CIPHERTEXT_WIDTH'd15473483;
publickey_row[5900] = `CIPHERTEXT_WIDTH'd1556195;
publickey_row[5901] = `CIPHERTEXT_WIDTH'd12370879;
publickey_row[5902] = `CIPHERTEXT_WIDTH'd4695233;
publickey_row[5903] = `CIPHERTEXT_WIDTH'd7449750;
publickey_row[5904] = `CIPHERTEXT_WIDTH'd15655847;
publickey_row[5905] = `CIPHERTEXT_WIDTH'd8414252;
publickey_row[5906] = `CIPHERTEXT_WIDTH'd2818945;
publickey_row[5907] = `CIPHERTEXT_WIDTH'd6685272;
publickey_row[5908] = `CIPHERTEXT_WIDTH'd15738641;
publickey_row[5909] = `CIPHERTEXT_WIDTH'd9030536;
publickey_row[5910] = `CIPHERTEXT_WIDTH'd12658037;
publickey_row[5911] = `CIPHERTEXT_WIDTH'd9520150;
publickey_row[5912] = `CIPHERTEXT_WIDTH'd15475527;
publickey_row[5913] = `CIPHERTEXT_WIDTH'd14596984;
publickey_row[5914] = `CIPHERTEXT_WIDTH'd825124;
publickey_row[5915] = `CIPHERTEXT_WIDTH'd3730202;
publickey_row[5916] = `CIPHERTEXT_WIDTH'd12825853;
publickey_row[5917] = `CIPHERTEXT_WIDTH'd16084139;
publickey_row[5918] = `CIPHERTEXT_WIDTH'd1462787;
publickey_row[5919] = `CIPHERTEXT_WIDTH'd4359983;
publickey_row[5920] = `CIPHERTEXT_WIDTH'd10106381;
publickey_row[5921] = `CIPHERTEXT_WIDTH'd2098594;
publickey_row[5922] = `CIPHERTEXT_WIDTH'd3949863;
publickey_row[5923] = `CIPHERTEXT_WIDTH'd1393852;
publickey_row[5924] = `CIPHERTEXT_WIDTH'd7939674;
publickey_row[5925] = `CIPHERTEXT_WIDTH'd4171657;
publickey_row[5926] = `CIPHERTEXT_WIDTH'd6137483;
publickey_row[5927] = `CIPHERTEXT_WIDTH'd8897975;
publickey_row[5928] = `CIPHERTEXT_WIDTH'd2836667;
publickey_row[5929] = `CIPHERTEXT_WIDTH'd5851305;
publickey_row[5930] = `CIPHERTEXT_WIDTH'd14518420;
publickey_row[5931] = `CIPHERTEXT_WIDTH'd4476115;
publickey_row[5932] = `CIPHERTEXT_WIDTH'd13281947;
publickey_row[5933] = `CIPHERTEXT_WIDTH'd3109461;
publickey_row[5934] = `CIPHERTEXT_WIDTH'd696246;
publickey_row[5935] = `CIPHERTEXT_WIDTH'd3865550;
publickey_row[5936] = `CIPHERTEXT_WIDTH'd5912885;
publickey_row[5937] = `CIPHERTEXT_WIDTH'd5390895;
publickey_row[5938] = `CIPHERTEXT_WIDTH'd11423884;
publickey_row[5939] = `CIPHERTEXT_WIDTH'd10498249;
publickey_row[5940] = `CIPHERTEXT_WIDTH'd3274738;
publickey_row[5941] = `CIPHERTEXT_WIDTH'd5977249;
publickey_row[5942] = `CIPHERTEXT_WIDTH'd16178189;
publickey_row[5943] = `CIPHERTEXT_WIDTH'd6570312;
publickey_row[5944] = `CIPHERTEXT_WIDTH'd4941115;
publickey_row[5945] = `CIPHERTEXT_WIDTH'd9959168;
publickey_row[5946] = `CIPHERTEXT_WIDTH'd12351582;
publickey_row[5947] = `CIPHERTEXT_WIDTH'd11915486;
publickey_row[5948] = `CIPHERTEXT_WIDTH'd10995859;
publickey_row[5949] = `CIPHERTEXT_WIDTH'd16008433;
publickey_row[5950] = `CIPHERTEXT_WIDTH'd14242627;
publickey_row[5951] = `CIPHERTEXT_WIDTH'd16320055;
publickey_row[5952] = `CIPHERTEXT_WIDTH'd1623508;
publickey_row[5953] = `CIPHERTEXT_WIDTH'd4870078;
publickey_row[5954] = `CIPHERTEXT_WIDTH'd5203366;
publickey_row[5955] = `CIPHERTEXT_WIDTH'd8163579;
publickey_row[5956] = `CIPHERTEXT_WIDTH'd12040571;
publickey_row[5957] = `CIPHERTEXT_WIDTH'd15908412;
publickey_row[5958] = `CIPHERTEXT_WIDTH'd9835235;
publickey_row[5959] = `CIPHERTEXT_WIDTH'd7294060;
publickey_row[5960] = `CIPHERTEXT_WIDTH'd12287935;
publickey_row[5961] = `CIPHERTEXT_WIDTH'd12612665;
publickey_row[5962] = `CIPHERTEXT_WIDTH'd3462481;
publickey_row[5963] = `CIPHERTEXT_WIDTH'd9526877;
publickey_row[5964] = `CIPHERTEXT_WIDTH'd15935268;
publickey_row[5965] = `CIPHERTEXT_WIDTH'd1434735;
publickey_row[5966] = `CIPHERTEXT_WIDTH'd2082015;
publickey_row[5967] = `CIPHERTEXT_WIDTH'd9115598;
publickey_row[5968] = `CIPHERTEXT_WIDTH'd3589178;
publickey_row[5969] = `CIPHERTEXT_WIDTH'd16043672;
publickey_row[5970] = `CIPHERTEXT_WIDTH'd13045664;
publickey_row[5971] = `CIPHERTEXT_WIDTH'd10628404;
publickey_row[5972] = `CIPHERTEXT_WIDTH'd984621;
publickey_row[5973] = `CIPHERTEXT_WIDTH'd2724577;
publickey_row[5974] = `CIPHERTEXT_WIDTH'd4740707;
publickey_row[5975] = `CIPHERTEXT_WIDTH'd6331592;
publickey_row[5976] = `CIPHERTEXT_WIDTH'd10883487;
publickey_row[5977] = `CIPHERTEXT_WIDTH'd4794510;
publickey_row[5978] = `CIPHERTEXT_WIDTH'd4281507;
publickey_row[5979] = `CIPHERTEXT_WIDTH'd12099165;
publickey_row[5980] = `CIPHERTEXT_WIDTH'd14511216;
publickey_row[5981] = `CIPHERTEXT_WIDTH'd6583309;
publickey_row[5982] = `CIPHERTEXT_WIDTH'd9620652;
publickey_row[5983] = `CIPHERTEXT_WIDTH'd13729750;
publickey_row[5984] = `CIPHERTEXT_WIDTH'd13719792;
publickey_row[5985] = `CIPHERTEXT_WIDTH'd10481654;
publickey_row[5986] = `CIPHERTEXT_WIDTH'd6727754;
publickey_row[5987] = `CIPHERTEXT_WIDTH'd15338955;
publickey_row[5988] = `CIPHERTEXT_WIDTH'd1295234;
publickey_row[5989] = `CIPHERTEXT_WIDTH'd6169374;
publickey_row[5990] = `CIPHERTEXT_WIDTH'd387016;
publickey_row[5991] = `CIPHERTEXT_WIDTH'd6893365;
publickey_row[5992] = `CIPHERTEXT_WIDTH'd16159208;
publickey_row[5993] = `CIPHERTEXT_WIDTH'd6775079;
publickey_row[5994] = `CIPHERTEXT_WIDTH'd5250689;
publickey_row[5995] = `CIPHERTEXT_WIDTH'd15738442;
publickey_row[5996] = `CIPHERTEXT_WIDTH'd7282324;
publickey_row[5997] = `CIPHERTEXT_WIDTH'd15563917;
publickey_row[5998] = `CIPHERTEXT_WIDTH'd4919231;
publickey_row[5999] = `CIPHERTEXT_WIDTH'd1402596;
publickey_row[6000] = `CIPHERTEXT_WIDTH'd14841621;
publickey_row[6001] = `CIPHERTEXT_WIDTH'd15027512;
publickey_row[6002] = `CIPHERTEXT_WIDTH'd5187138;
publickey_row[6003] = `CIPHERTEXT_WIDTH'd4943996;
publickey_row[6004] = `CIPHERTEXT_WIDTH'd13205828;
publickey_row[6005] = `CIPHERTEXT_WIDTH'd9974509;
publickey_row[6006] = `CIPHERTEXT_WIDTH'd12849083;
publickey_row[6007] = `CIPHERTEXT_WIDTH'd13391387;
publickey_row[6008] = `CIPHERTEXT_WIDTH'd10198640;
publickey_row[6009] = `CIPHERTEXT_WIDTH'd13279306;
publickey_row[6010] = `CIPHERTEXT_WIDTH'd15678936;
publickey_row[6011] = `CIPHERTEXT_WIDTH'd9224828;
publickey_row[6012] = `CIPHERTEXT_WIDTH'd8232513;
publickey_row[6013] = `CIPHERTEXT_WIDTH'd5371843;
publickey_row[6014] = `CIPHERTEXT_WIDTH'd13643563;
publickey_row[6015] = `CIPHERTEXT_WIDTH'd9352805;
publickey_row[6016] = `CIPHERTEXT_WIDTH'd12002774;
publickey_row[6017] = `CIPHERTEXT_WIDTH'd7280771;
publickey_row[6018] = `CIPHERTEXT_WIDTH'd13661904;
publickey_row[6019] = `CIPHERTEXT_WIDTH'd12906771;
publickey_row[6020] = `CIPHERTEXT_WIDTH'd6810299;
publickey_row[6021] = `CIPHERTEXT_WIDTH'd15987394;
publickey_row[6022] = `CIPHERTEXT_WIDTH'd3146492;
publickey_row[6023] = `CIPHERTEXT_WIDTH'd16498194;
publickey_row[6024] = `CIPHERTEXT_WIDTH'd6014632;
publickey_row[6025] = `CIPHERTEXT_WIDTH'd7867519;
publickey_row[6026] = `CIPHERTEXT_WIDTH'd5313609;
publickey_row[6027] = `CIPHERTEXT_WIDTH'd4788653;
publickey_row[6028] = `CIPHERTEXT_WIDTH'd5476287;
publickey_row[6029] = `CIPHERTEXT_WIDTH'd6983490;
publickey_row[6030] = `CIPHERTEXT_WIDTH'd1287088;
publickey_row[6031] = `CIPHERTEXT_WIDTH'd7330505;
publickey_row[6032] = `CIPHERTEXT_WIDTH'd2062037;
publickey_row[6033] = `CIPHERTEXT_WIDTH'd5240421;
publickey_row[6034] = `CIPHERTEXT_WIDTH'd5676809;
publickey_row[6035] = `CIPHERTEXT_WIDTH'd1388777;
publickey_row[6036] = `CIPHERTEXT_WIDTH'd15284567;
publickey_row[6037] = `CIPHERTEXT_WIDTH'd6653571;
publickey_row[6038] = `CIPHERTEXT_WIDTH'd14951922;
publickey_row[6039] = `CIPHERTEXT_WIDTH'd14190163;
publickey_row[6040] = `CIPHERTEXT_WIDTH'd16090822;
publickey_row[6041] = `CIPHERTEXT_WIDTH'd9690032;
publickey_row[6042] = `CIPHERTEXT_WIDTH'd11926378;
publickey_row[6043] = `CIPHERTEXT_WIDTH'd15779077;
publickey_row[6044] = `CIPHERTEXT_WIDTH'd7406336;
publickey_row[6045] = `CIPHERTEXT_WIDTH'd13362847;
publickey_row[6046] = `CIPHERTEXT_WIDTH'd8672906;
publickey_row[6047] = `CIPHERTEXT_WIDTH'd5699438;
publickey_row[6048] = `CIPHERTEXT_WIDTH'd6855401;
publickey_row[6049] = `CIPHERTEXT_WIDTH'd1426453;
publickey_row[6050] = `CIPHERTEXT_WIDTH'd3453738;
publickey_row[6051] = `CIPHERTEXT_WIDTH'd15949384;
publickey_row[6052] = `CIPHERTEXT_WIDTH'd1435006;
publickey_row[6053] = `CIPHERTEXT_WIDTH'd9198355;
publickey_row[6054] = `CIPHERTEXT_WIDTH'd13021148;
publickey_row[6055] = `CIPHERTEXT_WIDTH'd7385150;
publickey_row[6056] = `CIPHERTEXT_WIDTH'd11857631;
publickey_row[6057] = `CIPHERTEXT_WIDTH'd11453957;
publickey_row[6058] = `CIPHERTEXT_WIDTH'd762958;
publickey_row[6059] = `CIPHERTEXT_WIDTH'd429742;
publickey_row[6060] = `CIPHERTEXT_WIDTH'd5318469;
publickey_row[6061] = `CIPHERTEXT_WIDTH'd12809696;
publickey_row[6062] = `CIPHERTEXT_WIDTH'd12072536;
publickey_row[6063] = `CIPHERTEXT_WIDTH'd10938591;
publickey_row[6064] = `CIPHERTEXT_WIDTH'd7440347;
publickey_row[6065] = `CIPHERTEXT_WIDTH'd13341630;
publickey_row[6066] = `CIPHERTEXT_WIDTH'd10478174;
publickey_row[6067] = `CIPHERTEXT_WIDTH'd15185281;
publickey_row[6068] = `CIPHERTEXT_WIDTH'd9929221;
publickey_row[6069] = `CIPHERTEXT_WIDTH'd13234728;
publickey_row[6070] = `CIPHERTEXT_WIDTH'd14811872;
publickey_row[6071] = `CIPHERTEXT_WIDTH'd13843548;
publickey_row[6072] = `CIPHERTEXT_WIDTH'd16293455;
publickey_row[6073] = `CIPHERTEXT_WIDTH'd7115318;
publickey_row[6074] = `CIPHERTEXT_WIDTH'd11541245;
publickey_row[6075] = `CIPHERTEXT_WIDTH'd4706168;
publickey_row[6076] = `CIPHERTEXT_WIDTH'd7475814;
publickey_row[6077] = `CIPHERTEXT_WIDTH'd6926916;
publickey_row[6078] = `CIPHERTEXT_WIDTH'd5242087;
publickey_row[6079] = `CIPHERTEXT_WIDTH'd15959335;
publickey_row[6080] = `CIPHERTEXT_WIDTH'd4949740;
publickey_row[6081] = `CIPHERTEXT_WIDTH'd8996465;
publickey_row[6082] = `CIPHERTEXT_WIDTH'd3106676;
publickey_row[6083] = `CIPHERTEXT_WIDTH'd10167571;
publickey_row[6084] = `CIPHERTEXT_WIDTH'd5097501;
publickey_row[6085] = `CIPHERTEXT_WIDTH'd15054730;
publickey_row[6086] = `CIPHERTEXT_WIDTH'd5881643;
publickey_row[6087] = `CIPHERTEXT_WIDTH'd10022124;
publickey_row[6088] = `CIPHERTEXT_WIDTH'd10905975;
publickey_row[6089] = `CIPHERTEXT_WIDTH'd2050624;
publickey_row[6090] = `CIPHERTEXT_WIDTH'd12052149;
publickey_row[6091] = `CIPHERTEXT_WIDTH'd14067300;
publickey_row[6092] = `CIPHERTEXT_WIDTH'd10675153;
publickey_row[6093] = `CIPHERTEXT_WIDTH'd200620;
publickey_row[6094] = `CIPHERTEXT_WIDTH'd2819550;
publickey_row[6095] = `CIPHERTEXT_WIDTH'd7714523;
publickey_row[6096] = `CIPHERTEXT_WIDTH'd10882802;
publickey_row[6097] = `CIPHERTEXT_WIDTH'd15143056;
publickey_row[6098] = `CIPHERTEXT_WIDTH'd11728061;
publickey_row[6099] = `CIPHERTEXT_WIDTH'd6737120;
publickey_row[6100] = `CIPHERTEXT_WIDTH'd1433455;
publickey_row[6101] = `CIPHERTEXT_WIDTH'd14041316;
publickey_row[6102] = `CIPHERTEXT_WIDTH'd4532273;
publickey_row[6103] = `CIPHERTEXT_WIDTH'd9851556;
publickey_row[6104] = `CIPHERTEXT_WIDTH'd1108000;
publickey_row[6105] = `CIPHERTEXT_WIDTH'd13747802;
publickey_row[6106] = `CIPHERTEXT_WIDTH'd7415441;
publickey_row[6107] = `CIPHERTEXT_WIDTH'd13522710;
publickey_row[6108] = `CIPHERTEXT_WIDTH'd1546107;
publickey_row[6109] = `CIPHERTEXT_WIDTH'd2733758;
publickey_row[6110] = `CIPHERTEXT_WIDTH'd5048322;
publickey_row[6111] = `CIPHERTEXT_WIDTH'd9144289;
publickey_row[6112] = `CIPHERTEXT_WIDTH'd3477120;
publickey_row[6113] = `CIPHERTEXT_WIDTH'd10877561;
publickey_row[6114] = `CIPHERTEXT_WIDTH'd13435839;
publickey_row[6115] = `CIPHERTEXT_WIDTH'd14930676;
publickey_row[6116] = `CIPHERTEXT_WIDTH'd2385798;
publickey_row[6117] = `CIPHERTEXT_WIDTH'd5904826;
publickey_row[6118] = `CIPHERTEXT_WIDTH'd2605868;
publickey_row[6119] = `CIPHERTEXT_WIDTH'd10958022;
publickey_row[6120] = `CIPHERTEXT_WIDTH'd11636151;
publickey_row[6121] = `CIPHERTEXT_WIDTH'd768826;
publickey_row[6122] = `CIPHERTEXT_WIDTH'd13293599;
publickey_row[6123] = `CIPHERTEXT_WIDTH'd1819387;
publickey_row[6124] = `CIPHERTEXT_WIDTH'd3508070;
publickey_row[6125] = `CIPHERTEXT_WIDTH'd15330840;
publickey_row[6126] = `CIPHERTEXT_WIDTH'd4636605;
publickey_row[6127] = `CIPHERTEXT_WIDTH'd9696619;
publickey_row[6128] = `CIPHERTEXT_WIDTH'd12427809;
publickey_row[6129] = `CIPHERTEXT_WIDTH'd4636615;
publickey_row[6130] = `CIPHERTEXT_WIDTH'd4934083;
publickey_row[6131] = `CIPHERTEXT_WIDTH'd12093174;
publickey_row[6132] = `CIPHERTEXT_WIDTH'd6537204;
publickey_row[6133] = `CIPHERTEXT_WIDTH'd12100956;
publickey_row[6134] = `CIPHERTEXT_WIDTH'd9742450;
publickey_row[6135] = `CIPHERTEXT_WIDTH'd1120219;
publickey_row[6136] = `CIPHERTEXT_WIDTH'd15633979;
publickey_row[6137] = `CIPHERTEXT_WIDTH'd683645;
publickey_row[6138] = `CIPHERTEXT_WIDTH'd8940450;
publickey_row[6139] = `CIPHERTEXT_WIDTH'd16106124;
publickey_row[6140] = `CIPHERTEXT_WIDTH'd997679;
publickey_row[6141] = `CIPHERTEXT_WIDTH'd16448367;
publickey_row[6142] = `CIPHERTEXT_WIDTH'd14534015;
publickey_row[6143] = `CIPHERTEXT_WIDTH'd3614139;
publickey_row[6144] = `CIPHERTEXT_WIDTH'd16602904;
publickey_row[6145] = `CIPHERTEXT_WIDTH'd16728028;
publickey_row[6146] = `CIPHERTEXT_WIDTH'd5868186;
publickey_row[6147] = `CIPHERTEXT_WIDTH'd1652096;
publickey_row[6148] = `CIPHERTEXT_WIDTH'd7498293;
publickey_row[6149] = `CIPHERTEXT_WIDTH'd11343085;
publickey_row[6150] = `CIPHERTEXT_WIDTH'd4073275;
publickey_row[6151] = `CIPHERTEXT_WIDTH'd2392849;
publickey_row[6152] = `CIPHERTEXT_WIDTH'd15392664;
publickey_row[6153] = `CIPHERTEXT_WIDTH'd11754556;
publickey_row[6154] = `CIPHERTEXT_WIDTH'd9180538;
publickey_row[6155] = `CIPHERTEXT_WIDTH'd5296949;
publickey_row[6156] = `CIPHERTEXT_WIDTH'd6159987;
publickey_row[6157] = `CIPHERTEXT_WIDTH'd14477686;
publickey_row[6158] = `CIPHERTEXT_WIDTH'd9711390;
publickey_row[6159] = `CIPHERTEXT_WIDTH'd14637832;
publickey_row[6160] = `CIPHERTEXT_WIDTH'd125191;
publickey_row[6161] = `CIPHERTEXT_WIDTH'd7305538;
publickey_row[6162] = `CIPHERTEXT_WIDTH'd14929737;
publickey_row[6163] = `CIPHERTEXT_WIDTH'd13543225;
publickey_row[6164] = `CIPHERTEXT_WIDTH'd3038054;
publickey_row[6165] = `CIPHERTEXT_WIDTH'd15413235;
publickey_row[6166] = `CIPHERTEXT_WIDTH'd374707;
publickey_row[6167] = `CIPHERTEXT_WIDTH'd11600140;
publickey_row[6168] = `CIPHERTEXT_WIDTH'd2474225;
publickey_row[6169] = `CIPHERTEXT_WIDTH'd3785245;
publickey_row[6170] = `CIPHERTEXT_WIDTH'd12642453;
publickey_row[6171] = `CIPHERTEXT_WIDTH'd4424274;
publickey_row[6172] = `CIPHERTEXT_WIDTH'd4034562;
publickey_row[6173] = `CIPHERTEXT_WIDTH'd13499427;
publickey_row[6174] = `CIPHERTEXT_WIDTH'd8190419;
publickey_row[6175] = `CIPHERTEXT_WIDTH'd7797442;
publickey_row[6176] = `CIPHERTEXT_WIDTH'd1381205;
publickey_row[6177] = `CIPHERTEXT_WIDTH'd8260858;
publickey_row[6178] = `CIPHERTEXT_WIDTH'd1790246;
publickey_row[6179] = `CIPHERTEXT_WIDTH'd14143447;
publickey_row[6180] = `CIPHERTEXT_WIDTH'd2708901;
publickey_row[6181] = `CIPHERTEXT_WIDTH'd3750287;
publickey_row[6182] = `CIPHERTEXT_WIDTH'd15133455;
publickey_row[6183] = `CIPHERTEXT_WIDTH'd5318521;
publickey_row[6184] = `CIPHERTEXT_WIDTH'd15051189;
publickey_row[6185] = `CIPHERTEXT_WIDTH'd10132493;
publickey_row[6186] = `CIPHERTEXT_WIDTH'd16342553;
publickey_row[6187] = `CIPHERTEXT_WIDTH'd15509061;
publickey_row[6188] = `CIPHERTEXT_WIDTH'd7934721;
publickey_row[6189] = `CIPHERTEXT_WIDTH'd380218;
publickey_row[6190] = `CIPHERTEXT_WIDTH'd4969920;
publickey_row[6191] = `CIPHERTEXT_WIDTH'd13970035;
publickey_row[6192] = `CIPHERTEXT_WIDTH'd12832969;
publickey_row[6193] = `CIPHERTEXT_WIDTH'd5902434;
publickey_row[6194] = `CIPHERTEXT_WIDTH'd93466;
publickey_row[6195] = `CIPHERTEXT_WIDTH'd3125701;
publickey_row[6196] = `CIPHERTEXT_WIDTH'd6416906;
publickey_row[6197] = `CIPHERTEXT_WIDTH'd8349007;
publickey_row[6198] = `CIPHERTEXT_WIDTH'd9126771;
publickey_row[6199] = `CIPHERTEXT_WIDTH'd6547358;
publickey_row[6200] = `CIPHERTEXT_WIDTH'd13457611;
publickey_row[6201] = `CIPHERTEXT_WIDTH'd11110402;
publickey_row[6202] = `CIPHERTEXT_WIDTH'd11396926;
publickey_row[6203] = `CIPHERTEXT_WIDTH'd10360847;
publickey_row[6204] = `CIPHERTEXT_WIDTH'd4321302;
publickey_row[6205] = `CIPHERTEXT_WIDTH'd9243445;
publickey_row[6206] = `CIPHERTEXT_WIDTH'd3254945;
publickey_row[6207] = `CIPHERTEXT_WIDTH'd12263113;
publickey_row[6208] = `CIPHERTEXT_WIDTH'd8223475;
publickey_row[6209] = `CIPHERTEXT_WIDTH'd6933141;
publickey_row[6210] = `CIPHERTEXT_WIDTH'd8631748;
publickey_row[6211] = `CIPHERTEXT_WIDTH'd3565507;
publickey_row[6212] = `CIPHERTEXT_WIDTH'd4542894;
publickey_row[6213] = `CIPHERTEXT_WIDTH'd6187005;
publickey_row[6214] = `CIPHERTEXT_WIDTH'd14750139;
publickey_row[6215] = `CIPHERTEXT_WIDTH'd1107786;
publickey_row[6216] = `CIPHERTEXT_WIDTH'd2014896;
publickey_row[6217] = `CIPHERTEXT_WIDTH'd5827636;
publickey_row[6218] = `CIPHERTEXT_WIDTH'd15033633;
publickey_row[6219] = `CIPHERTEXT_WIDTH'd16627078;
publickey_row[6220] = `CIPHERTEXT_WIDTH'd5099911;
publickey_row[6221] = `CIPHERTEXT_WIDTH'd10218896;
publickey_row[6222] = `CIPHERTEXT_WIDTH'd4455200;
publickey_row[6223] = `CIPHERTEXT_WIDTH'd10708116;
publickey_row[6224] = `CIPHERTEXT_WIDTH'd9584731;
publickey_row[6225] = `CIPHERTEXT_WIDTH'd8099147;
publickey_row[6226] = `CIPHERTEXT_WIDTH'd13756370;
publickey_row[6227] = `CIPHERTEXT_WIDTH'd13511891;
publickey_row[6228] = `CIPHERTEXT_WIDTH'd2019171;
publickey_row[6229] = `CIPHERTEXT_WIDTH'd8676508;
publickey_row[6230] = `CIPHERTEXT_WIDTH'd14698008;
publickey_row[6231] = `CIPHERTEXT_WIDTH'd7338681;
publickey_row[6232] = `CIPHERTEXT_WIDTH'd1287165;
publickey_row[6233] = `CIPHERTEXT_WIDTH'd12435404;
publickey_row[6234] = `CIPHERTEXT_WIDTH'd11487378;
publickey_row[6235] = `CIPHERTEXT_WIDTH'd3319659;
publickey_row[6236] = `CIPHERTEXT_WIDTH'd2514204;
publickey_row[6237] = `CIPHERTEXT_WIDTH'd16285099;
publickey_row[6238] = `CIPHERTEXT_WIDTH'd13233383;
publickey_row[6239] = `CIPHERTEXT_WIDTH'd14768493;
publickey_row[6240] = `CIPHERTEXT_WIDTH'd904908;
publickey_row[6241] = `CIPHERTEXT_WIDTH'd13262458;
publickey_row[6242] = `CIPHERTEXT_WIDTH'd9149106;
publickey_row[6243] = `CIPHERTEXT_WIDTH'd11837127;
publickey_row[6244] = `CIPHERTEXT_WIDTH'd1225838;
publickey_row[6245] = `CIPHERTEXT_WIDTH'd11764717;
publickey_row[6246] = `CIPHERTEXT_WIDTH'd12885625;
publickey_row[6247] = `CIPHERTEXT_WIDTH'd7425424;
publickey_row[6248] = `CIPHERTEXT_WIDTH'd7590961;
publickey_row[6249] = `CIPHERTEXT_WIDTH'd4440277;
publickey_row[6250] = `CIPHERTEXT_WIDTH'd3059080;
publickey_row[6251] = `CIPHERTEXT_WIDTH'd14341770;
publickey_row[6252] = `CIPHERTEXT_WIDTH'd10274922;
publickey_row[6253] = `CIPHERTEXT_WIDTH'd9741583;
publickey_row[6254] = `CIPHERTEXT_WIDTH'd4047273;
publickey_row[6255] = `CIPHERTEXT_WIDTH'd1085544;
publickey_row[6256] = `CIPHERTEXT_WIDTH'd10023805;
publickey_row[6257] = `CIPHERTEXT_WIDTH'd262704;
publickey_row[6258] = `CIPHERTEXT_WIDTH'd8184011;
publickey_row[6259] = `CIPHERTEXT_WIDTH'd6215723;
publickey_row[6260] = `CIPHERTEXT_WIDTH'd4273708;
publickey_row[6261] = `CIPHERTEXT_WIDTH'd8902061;
publickey_row[6262] = `CIPHERTEXT_WIDTH'd183469;
publickey_row[6263] = `CIPHERTEXT_WIDTH'd10165706;
publickey_row[6264] = `CIPHERTEXT_WIDTH'd5472778;
publickey_row[6265] = `CIPHERTEXT_WIDTH'd2581624;
publickey_row[6266] = `CIPHERTEXT_WIDTH'd5395529;
publickey_row[6267] = `CIPHERTEXT_WIDTH'd14979812;
publickey_row[6268] = `CIPHERTEXT_WIDTH'd11557804;
publickey_row[6269] = `CIPHERTEXT_WIDTH'd4719146;
publickey_row[6270] = `CIPHERTEXT_WIDTH'd16580087;
publickey_row[6271] = `CIPHERTEXT_WIDTH'd2792636;
publickey_row[6272] = `CIPHERTEXT_WIDTH'd8707829;
publickey_row[6273] = `CIPHERTEXT_WIDTH'd4548345;
publickey_row[6274] = `CIPHERTEXT_WIDTH'd6599347;
publickey_row[6275] = `CIPHERTEXT_WIDTH'd6933927;
publickey_row[6276] = `CIPHERTEXT_WIDTH'd6649663;
publickey_row[6277] = `CIPHERTEXT_WIDTH'd14258198;
publickey_row[6278] = `CIPHERTEXT_WIDTH'd11349601;
publickey_row[6279] = `CIPHERTEXT_WIDTH'd12169728;
publickey_row[6280] = `CIPHERTEXT_WIDTH'd14517097;
publickey_row[6281] = `CIPHERTEXT_WIDTH'd2565373;
publickey_row[6282] = `CIPHERTEXT_WIDTH'd11951073;
publickey_row[6283] = `CIPHERTEXT_WIDTH'd4171982;
publickey_row[6284] = `CIPHERTEXT_WIDTH'd3398328;
publickey_row[6285] = `CIPHERTEXT_WIDTH'd2610616;
publickey_row[6286] = `CIPHERTEXT_WIDTH'd9069320;
publickey_row[6287] = `CIPHERTEXT_WIDTH'd2845244;
publickey_row[6288] = `CIPHERTEXT_WIDTH'd1436132;
publickey_row[6289] = `CIPHERTEXT_WIDTH'd9472956;
publickey_row[6290] = `CIPHERTEXT_WIDTH'd12019127;
publickey_row[6291] = `CIPHERTEXT_WIDTH'd6055496;
publickey_row[6292] = `CIPHERTEXT_WIDTH'd13385173;
publickey_row[6293] = `CIPHERTEXT_WIDTH'd3374505;
publickey_row[6294] = `CIPHERTEXT_WIDTH'd13479244;
publickey_row[6295] = `CIPHERTEXT_WIDTH'd4553626;
publickey_row[6296] = `CIPHERTEXT_WIDTH'd13293572;
publickey_row[6297] = `CIPHERTEXT_WIDTH'd16219895;
publickey_row[6298] = `CIPHERTEXT_WIDTH'd6076313;
publickey_row[6299] = `CIPHERTEXT_WIDTH'd15924570;
publickey_row[6300] = `CIPHERTEXT_WIDTH'd12134916;
publickey_row[6301] = `CIPHERTEXT_WIDTH'd7162304;
publickey_row[6302] = `CIPHERTEXT_WIDTH'd15858856;
publickey_row[6303] = `CIPHERTEXT_WIDTH'd16553174;
publickey_row[6304] = `CIPHERTEXT_WIDTH'd16369960;
publickey_row[6305] = `CIPHERTEXT_WIDTH'd7092313;
publickey_row[6306] = `CIPHERTEXT_WIDTH'd4362559;
publickey_row[6307] = `CIPHERTEXT_WIDTH'd14545983;
publickey_row[6308] = `CIPHERTEXT_WIDTH'd13040984;
publickey_row[6309] = `CIPHERTEXT_WIDTH'd5883100;
publickey_row[6310] = `CIPHERTEXT_WIDTH'd15566451;
publickey_row[6311] = `CIPHERTEXT_WIDTH'd6267735;
publickey_row[6312] = `CIPHERTEXT_WIDTH'd13233157;
publickey_row[6313] = `CIPHERTEXT_WIDTH'd12933947;
publickey_row[6314] = `CIPHERTEXT_WIDTH'd92699;
publickey_row[6315] = `CIPHERTEXT_WIDTH'd1529015;
publickey_row[6316] = `CIPHERTEXT_WIDTH'd9054660;
publickey_row[6317] = `CIPHERTEXT_WIDTH'd10398230;
publickey_row[6318] = `CIPHERTEXT_WIDTH'd9252303;
publickey_row[6319] = `CIPHERTEXT_WIDTH'd978574;
publickey_row[6320] = `CIPHERTEXT_WIDTH'd13881858;
publickey_row[6321] = `CIPHERTEXT_WIDTH'd7034632;
publickey_row[6322] = `CIPHERTEXT_WIDTH'd1771111;
publickey_row[6323] = `CIPHERTEXT_WIDTH'd753407;
publickey_row[6324] = `CIPHERTEXT_WIDTH'd2458450;
publickey_row[6325] = `CIPHERTEXT_WIDTH'd15649597;
publickey_row[6326] = `CIPHERTEXT_WIDTH'd736838;
publickey_row[6327] = `CIPHERTEXT_WIDTH'd14463781;
publickey_row[6328] = `CIPHERTEXT_WIDTH'd13936670;
publickey_row[6329] = `CIPHERTEXT_WIDTH'd15881910;
publickey_row[6330] = `CIPHERTEXT_WIDTH'd9321147;
publickey_row[6331] = `CIPHERTEXT_WIDTH'd11021405;
publickey_row[6332] = `CIPHERTEXT_WIDTH'd3423997;
publickey_row[6333] = `CIPHERTEXT_WIDTH'd12858236;
publickey_row[6334] = `CIPHERTEXT_WIDTH'd4395062;
publickey_row[6335] = `CIPHERTEXT_WIDTH'd2919352;
publickey_row[6336] = `CIPHERTEXT_WIDTH'd13724740;
publickey_row[6337] = `CIPHERTEXT_WIDTH'd8599255;
publickey_row[6338] = `CIPHERTEXT_WIDTH'd7630065;
publickey_row[6339] = `CIPHERTEXT_WIDTH'd14680831;
publickey_row[6340] = `CIPHERTEXT_WIDTH'd12881767;
publickey_row[6341] = `CIPHERTEXT_WIDTH'd1973404;
publickey_row[6342] = `CIPHERTEXT_WIDTH'd14830325;
publickey_row[6343] = `CIPHERTEXT_WIDTH'd10800901;
publickey_row[6344] = `CIPHERTEXT_WIDTH'd8255020;
publickey_row[6345] = `CIPHERTEXT_WIDTH'd14110516;
publickey_row[6346] = `CIPHERTEXT_WIDTH'd10985182;
publickey_row[6347] = `CIPHERTEXT_WIDTH'd8186115;
publickey_row[6348] = `CIPHERTEXT_WIDTH'd8426834;
publickey_row[6349] = `CIPHERTEXT_WIDTH'd4928358;
publickey_row[6350] = `CIPHERTEXT_WIDTH'd5211412;
publickey_row[6351] = `CIPHERTEXT_WIDTH'd6965071;
publickey_row[6352] = `CIPHERTEXT_WIDTH'd11696209;
publickey_row[6353] = `CIPHERTEXT_WIDTH'd14334190;
publickey_row[6354] = `CIPHERTEXT_WIDTH'd11046271;
publickey_row[6355] = `CIPHERTEXT_WIDTH'd492497;
publickey_row[6356] = `CIPHERTEXT_WIDTH'd8213549;
publickey_row[6357] = `CIPHERTEXT_WIDTH'd5065159;
publickey_row[6358] = `CIPHERTEXT_WIDTH'd14215547;
publickey_row[6359] = `CIPHERTEXT_WIDTH'd7690610;
publickey_row[6360] = `CIPHERTEXT_WIDTH'd1080173;
publickey_row[6361] = `CIPHERTEXT_WIDTH'd15298258;
publickey_row[6362] = `CIPHERTEXT_WIDTH'd1318601;
publickey_row[6363] = `CIPHERTEXT_WIDTH'd1570810;
publickey_row[6364] = `CIPHERTEXT_WIDTH'd3447324;
publickey_row[6365] = `CIPHERTEXT_WIDTH'd7510262;
publickey_row[6366] = `CIPHERTEXT_WIDTH'd9719572;
publickey_row[6367] = `CIPHERTEXT_WIDTH'd10341779;
publickey_row[6368] = `CIPHERTEXT_WIDTH'd12768324;
publickey_row[6369] = `CIPHERTEXT_WIDTH'd6494200;
publickey_row[6370] = `CIPHERTEXT_WIDTH'd10626620;
publickey_row[6371] = `CIPHERTEXT_WIDTH'd10808382;
publickey_row[6372] = `CIPHERTEXT_WIDTH'd447211;
publickey_row[6373] = `CIPHERTEXT_WIDTH'd8252186;
publickey_row[6374] = `CIPHERTEXT_WIDTH'd15609984;
publickey_row[6375] = `CIPHERTEXT_WIDTH'd7737098;
publickey_row[6376] = `CIPHERTEXT_WIDTH'd13575139;
publickey_row[6377] = `CIPHERTEXT_WIDTH'd16331366;
publickey_row[6378] = `CIPHERTEXT_WIDTH'd14576780;
publickey_row[6379] = `CIPHERTEXT_WIDTH'd7329576;
publickey_row[6380] = `CIPHERTEXT_WIDTH'd1740604;
publickey_row[6381] = `CIPHERTEXT_WIDTH'd5073721;
publickey_row[6382] = `CIPHERTEXT_WIDTH'd4932276;
publickey_row[6383] = `CIPHERTEXT_WIDTH'd13485836;
publickey_row[6384] = `CIPHERTEXT_WIDTH'd10936537;
publickey_row[6385] = `CIPHERTEXT_WIDTH'd11869276;
publickey_row[6386] = `CIPHERTEXT_WIDTH'd12373621;
publickey_row[6387] = `CIPHERTEXT_WIDTH'd6304954;
publickey_row[6388] = `CIPHERTEXT_WIDTH'd15476159;
publickey_row[6389] = `CIPHERTEXT_WIDTH'd14576791;
publickey_row[6390] = `CIPHERTEXT_WIDTH'd9409456;
publickey_row[6391] = `CIPHERTEXT_WIDTH'd9941786;
publickey_row[6392] = `CIPHERTEXT_WIDTH'd5154441;
publickey_row[6393] = `CIPHERTEXT_WIDTH'd4963868;
publickey_row[6394] = `CIPHERTEXT_WIDTH'd1122045;
publickey_row[6395] = `CIPHERTEXT_WIDTH'd11880790;
publickey_row[6396] = `CIPHERTEXT_WIDTH'd16657171;
publickey_row[6397] = `CIPHERTEXT_WIDTH'd11665055;
publickey_row[6398] = `CIPHERTEXT_WIDTH'd8322935;
publickey_row[6399] = `CIPHERTEXT_WIDTH'd8002302;
publickey_row[6400] = `CIPHERTEXT_WIDTH'd674431;
publickey_row[6401] = `CIPHERTEXT_WIDTH'd16751942;
publickey_row[6402] = `CIPHERTEXT_WIDTH'd6000123;
publickey_row[6403] = `CIPHERTEXT_WIDTH'd5742877;
publickey_row[6404] = `CIPHERTEXT_WIDTH'd12960896;
publickey_row[6405] = `CIPHERTEXT_WIDTH'd10645910;
publickey_row[6406] = `CIPHERTEXT_WIDTH'd16037523;
publickey_row[6407] = `CIPHERTEXT_WIDTH'd9913274;
publickey_row[6408] = `CIPHERTEXT_WIDTH'd10681949;
publickey_row[6409] = `CIPHERTEXT_WIDTH'd7492691;
publickey_row[6410] = `CIPHERTEXT_WIDTH'd5957866;
publickey_row[6411] = `CIPHERTEXT_WIDTH'd3126682;
publickey_row[6412] = `CIPHERTEXT_WIDTH'd1880436;
publickey_row[6413] = `CIPHERTEXT_WIDTH'd4451536;
publickey_row[6414] = `CIPHERTEXT_WIDTH'd12093192;
publickey_row[6415] = `CIPHERTEXT_WIDTH'd15973565;
publickey_row[6416] = `CIPHERTEXT_WIDTH'd1460509;
publickey_row[6417] = `CIPHERTEXT_WIDTH'd16450632;
publickey_row[6418] = `CIPHERTEXT_WIDTH'd12025906;
publickey_row[6419] = `CIPHERTEXT_WIDTH'd1566314;
publickey_row[6420] = `CIPHERTEXT_WIDTH'd8374026;
publickey_row[6421] = `CIPHERTEXT_WIDTH'd14891756;
publickey_row[6422] = `CIPHERTEXT_WIDTH'd13352027;
publickey_row[6423] = `CIPHERTEXT_WIDTH'd4409166;
publickey_row[6424] = `CIPHERTEXT_WIDTH'd7860522;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd0;
noise_select = `BIG_N'b00000110110111010010000101100111111100101001100111001101110011110110101111010111101010010110000001111110111100011010011110000001101001010110001110110101100100110000110100011111011100000100111101010011011011110001001011010010001111011100011010010101010110100001001101101010000111001000010101101100101100100110110010000000111100001100100110100001111100000110111010110100011100101001010101101101100000000000110100110101000101100101100010001101101010110111101001100100000000110100001001010011001001100001111111000110110111101101000000100011011000011111000010101000010011100110001001010110001110110011101010000011110110011011111001000001101100000100010101010010010111101010110010101101101011101001111001000110110110011001000010010011110010000110001101111011110011111010001110011110100111101110011011010111011001001000000111101111100001101001110000000110000010111000110101011010111100010011111000011101110101101001010000000001000100011001010001110111011001111101010001100011100011000011111010001100000110101000100011010010110101100111010010111101001000101101001010001111001010100100000001100000001101000010010011001000100000010000000101011011100000001010101001101111010101001100011010101011010110110110111011000111001000101011010001101010000100101001001001100011010100101110010000100000101100000001101011001010110111011011100101000001111000000001110010001101111001111110110101101000100110101010010000111111000010010110000010101111001000011101001000011000100001101111111110110000111100001011001111000110000011011001001000000111111101110111011000010011000110000111000010001011010000110111011100000011100110110111110100010011100100000101000010001010001000110111100110011001000010001011110101111111111001111110111000000110110101011001001101100010101000010101101100100111100101011110000000001010101100100000010000101010000000010010011011001010011001001000110101011010001010110001111110110000100110111011111111110110110110111100111010000111111010001010011101010001110101000000101110000111100011011001101100000010000100110011000101110010001110111010010111101101110110010010110110100100110000011010001000111001111110111000011010011100101110000000000100010001110000110010110110100011011101111010011100000010000101101000010111100010010101111001001110111101001000100000101111111001001000110001001110011011010001000000101101101011101000011110000100011000111101110000001110111101101000111110100001001000111100100001010000101011011111111010100101000111110001101010110001110110001100010101000100110011000010010001100001000111111010000110001000110001111101100000100000110001110101111100110111010011000010010100100100111110110010101110110001011110111001111000101000001011100110111010000110000111111100110111011010100010010011011101111110100001100110001011011110011111011010001100111101111010001101000000101110101010000010101110100110010001100101111110011001011111111111000010100000000101011100100101111101011101101010111101011010100001000000010100000111110111101011101101000100011001110001010010001100011101010111001111100111000100001011110100011111001110110010111100000101111011110001000100000111110100110001100001101010101100110111110110101110011100011011000011011100010101010001001011011110101101000111010101010111111011011110000000100110101100011001100100110000101111110110001001100000010000010101101100001111000111000010010011110110111010101011000000111111111010010111000111111110101101001111101100000110000001100101001101101001000000001111100001110100100101111101010101000111010100100000001000001110000100010111010001101011101110011010100010001011011101101000000001101001101100011101000010110000000100110111110000011000010110011100101010111001011101001111100101111001111000001101010010101100011001100100010110110101010100101111001010100001101011100001010110000010100101101001010110101011001000001100011001010000100010000111100100001000000001101101100010111010001110011110010000110010010111110000110001110011101100001010110001110001101100001000110010110010001100100111101010001010000011010000000101111001111011010010010001101011101010101010100000110111110011001101010001011100101010110101001100010100001000110001000000110010001110110010000000011000010100000011101111000111011111010011010000001011010101111011010100011110110100000001010111111000110000100001010001111110100110111001001000000011010110101101001100111000011000001100000101011111000011101001001010000101000000101001110100011011100010011110000111100111011011110101111000110011001010101110010011111001110100010010111110101001100110010110010100000110000001011011111000101000011011100110111010010110110001001110000001100011010011110001100101111011100011001100100101010110110000100001101100110000001111000000011001100011010111101010000110010101011101001001101011000010111101110000010100010111110100100011010001100101111111001000100000000001010011111011000001011001000111001011010010011001011100100010011001101110111111101111001101100000110110010000011001111001001100100001000111100011111010110000111011101000001001111001101010011111101111011010010000011001011101010001000011101111100101101011101001110010010001010011010010100011111000000100110000111011110011001011101001011100010001111011100111100010010000011110001111001111110000101101101011100100111100101101110000001101000011101111000100110101101001100000011100110000111010100011111000000101000010001110110101011000010010101011100111011111001001110010011011100100101101110001010010101111101111000010110101100101110001011110101001000110000101001111100000010011111000111011101000000010101000110001011101010010110110100110101100001000101010111000110110100010101000111001100111000110101101111000110011011010011111111000111100011110011100001011011011010101011000001010011100111111110010110001001100100101010100111011001000101100101110011100001100100110000010011010000011001011011111010101111001100011010101000100110010111010010011010100010001010100001111111100111011000101111111111011010001101100010010111011011000110111111001001101110101011011101011110110000011100100011001010101110011010000010011010111100010101100110110000011000111000110111101110010010110011000011010101110110100001100110100011001011001101100101011000110101011010011100010011011101100000001111000100111111011101010111100000110111101001110101100100110001111101100001100010001010011100110111110011000011001001011111110010000000101110001100001100100011100011011101100011110000011111101001000110011011110001000101001001111100000011010101010100111110010010101101000110101010;
expected = 4685902;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);
#20;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd1;
noise_select = `BIG_N'b00011010011110100000110110001000000011001100011111111110001010110110001101101001000011000110111110110111101001010010100011010101001111010100001010000100000000110000011001000011100101000000110100010100000101010011100100111010110101110100101111000001100001111101000100101011001000010001100010111100110110001100000011001101000010101001100011000110011101010100000000111110101001100001011111101101110110000111000110000001100110100110011011111101011011110110010110100000000000101111010010101010011100110011111110010100010101010110001000111001101100000111011111000000000100011111000110101000001110100010001011000010110011010011000010111111111101101101000001100001010000000110001000110110000011100100010001111000100110000100111100111111001010100100010100011000111111001001100001010011100101101001000010000001111001101110100110010001110000010010100100110100101010100010000011001100101001100011011101110010000011110001000111000000001000000010011101001010010100001011001100100111100001101111111011111000011010011001011011111000101011111010110110110111011111011101011110000000111100011010001111001011001010000110111000010010000101110001111000011001001111011001010111100000110001111110101100110001001010001110110111001010000101001010001101100001100110011101001111000111110000010110111111011010101110000000111001110000111001101111100101000000011000101110011111101111011010001011101110010011001101110000001000010000100111100110010100101000111010111100111110100011001101010100001111000111010011100101000110010100011101000101100010011010000100001001111110011010001101111110111000000101110100101110110111010100000000110000110100000100111100110101101110111010100001011101001010011001011100101001101101010001110010110010011100111101010011101011111010100111011100100001000100000001011101011100000110110100111101101001011001110111010010001001101101011000000010001001100111101111000101111001000010111111001011111000011000001100111110010010111001100101100100101101101011011111000010010011010110101001101111100000100110111000011111101011000011101010010011100001000010111011111001110001010100010110100010101000110101101001100001010011111001011000011110011110101101011001100000010100101101111110101011101101100011000010011101000101010010011000100010000110001001010011101001100111100110111010100010000001010101011111110001101010011111010111011001110010001111101011010100101001100011111010000100010111111000111001111100110101111011110011111000001001100010111100000100100110110101111011101010100001000100100100000110000101101011011000100101011110010000001000010100100010111011000000010010011101101111101011101000000011000001111011100101011001010001001101010110001001111011001001110110100001000101001011001010000000111011001100011010001011001101010110011010111110010000010111111100000111010000100101101101001001101001011010110000111100110011111000011011000110110000111001110000001100110001111011011001000100000011100011111011010100000110100010010000111110110110010100100100100000101100100010110111100100110101001111100101010000011110000101111001001100111000111110011001001110111010010010001001101101111101101100101100111011100010100000001111100110110001011001001000000101110101000110001100100100001101010101010001000111000101101101101100111000001001111000000111011100000110101101001010011010110100010010000101010100010101000100101000000010110010001001100101100100111000000111010000110110010001011110010111100001010100011001010000001111111000110111101011100110001111111100110110101101010010000011011010111100000000110010011011101110000101010110111010011100111011101010111011100111000101110001000000001111101110001000100100011101111110111101100000011010101111000000001001000010011100010010010001010000101100000111001011001000011010001011101101010111001011001110010000111100101111000011011110101101100000110111101100000001000101100001010000110100000111011010111000110100111001110001001011001101100101011010110110001001011001011101101111110011111010000100110011111000010000110001001000100001100100110010111101001010010110001101001010010110010011011011110100101100101110110101011110011100001101010001111010001110101000100111001101001101001100101001011011001101111011001101000011011110011000000110001001101001101101100111011100100100000001101000000110100110111110100111110110101101000110111100110100000011001110110010111000000100101011110111111011111000001101100001100100101111010010101100111001011000001000000100001000111010001101001100111011111011010001101111101101111101010101010011100111110001001000101111010100001001100111011000001010110001101111110100100000100111111011000001100111111111010010110101000111111111001000111110000111101000010110110001111011000010100001000000110000000100110011000001000111001110001010000010000110000001011011000011111100011000010101000110010111010000111010110110100111010010110001011010111100011100111011111001101010111100001110101111011110110101100101010001100100101010010011001000100010111001110111111101111010010011000111000010100001111101101011010111111110000001010010111010000100110100000000001111101101110101010000111000000110010100001001111001101001111000011101100000111101000010000101000011110100101011010111010001000010011010101100011100111100101111100001010100011001010100100100110101010011000000001000001101101101110001011011001000011001000110101011110110111000111010111001010000110001101001011010001001011111111001001110111101111011010111111111000111010100101011010000010011010100000011110011110010111011110101001101001101110111011010111100110000111100011111101101011111110100111111100111101111100100110010111100010011110001010010110011011001101001100011000011101000001011111000111100111011100000110101110010011000001001110100001101010000111001010000000000101111110000000001111010010000101111111111011011000000110101011000010111110010110101001110111011000101011111001110100010000101111000001011100101100100101101101110111011101101001000011011001010110011000111100010110001101110011000001001101101001110011000111101100101101011110100010111110010001011010000111011001011011000111000001001011001101011011100000101001000101111001100001100001100110001000001110001101011010001110101100010110010100001011100110101101101111001100100001111111100110110100011100000110101110110101101000011001110101011010110111111000010011111100100101110010111100000100011110011110111110110000111101011001100000101000111101001001101001110011010110010110001101000101110101001000110100111011011010110100100000011011001110100000111101100100101000;
expected = 3580395;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);
#20;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd2;
noise_select = `BIG_N'b11101110110110001101100000111010000011101101110001101011010001000111100101010000011011000010110110001111100110010110000000100011000101000111000101111101000001101010001101101010011011110101000100010001100101001011100101111001001111101011001101110000110011101000010001010010011011100100100011011100110110101000000001100100100010110111010000001011101100100100110010110110101110100100101110111111011101000001110000111011010111100010101101011010111001001101110010100011101001101111100111010111001110011011100110010011011100101011010101101111010010110011001110000101100001001001101110101000101000111100010110100110010010000100011011010100111000000111100000100001010110010000000011010100110010101001001001101010110100100100010000011100111110011011111010000111001011100000110110100011110001100001110000011001101000010101001010010000000010001001010100001100001101000101010111100011101011001010011011001011110000101001001010010001111010000111110000001000001110101101000101010000010001001011011001100001001100100010101110101011001010101100010001000101000010100010001001000100010100110100101110101001101110000001111011111010011100111011011101010011011110101000010111011100001100001111111101010010010100101010011000010110100100101011111000000100100001000101100011010011111101101001011010100000001011101000000101001000100101001001011111110101110000111101101110000101000011000111101111010101000000101110111111110011101001010101110101000100011000010110010001000101011110101111011010001010011111101011101011101000101000010100010010010001110001101111010100011000100100001111000011000110010100101011100111110101001000011101001111010001110000001001010011110011011111101111101010001001101011010011001101101100011111100001111100010011110100110000110110001111000111110101100001111011000001010101111101111110000011111110011000010111101000101101001011000000000101110011011100001110000110011111001010111000100101010100011000010001001001110001000111011010011000111000110111000110111111011110011001001000101111011111111010101110011010111001111001000111111100110011001100110001011011001101000110111010000100101101011001110110111001101010010000001100100101011010001101101111110011001010101110001010011111101111001111001100101100101110110110001000011011011111000111100001010111111110110001010101100101001111011000101100000111000000110000110001110100100100101111010100100110000111100110101001000111110001100111000010011000111110101011010110010110100101111001101111011110000010001000101100101010100011111010001101111010111011011101000111001011110111110001111011011101000010100110000001101001100110111011001011011000011110100011000101000111111110101110010011110100000011110111000010001010100110101010011110110001010110111101000001000011010100010100110100110011000110010100000001001001101011011100000010110100001011000000010001101110100001010110011011011011110001110100000011010100101101010001110000000110111110001100111001010011000100000101000010000111010001110101111000110100001110101101100100110111011010101101110100110111110111010010101000000101001110101001000000100001110000011101100000110001110110011101011101110111101101111011101111101010010000011000111010100111110011000100101110101111101111011111101010010110101100111000110010001100100111010010001100111101110101001100010101010111100111111000011011101011101001111110111001010111111010101111110010100001001000010111110001110001110100111110001010110110110100111100111101110100100011000011001110100110110000010010101101111010110111000101001010100001100110111110100000111111101100100011011010110000011001110100110000100110100110001100100100011111010001111001111010100000100111000011111010111110010001011010001111011010001010000000101011100110001111110101101011110011000011101110100011010001000000000100010100000101111001001000111110100110101001001101101111011100010111110010001100110010010110101101110110001100011000111001010000010001101111100100001001111011001101011110111001010000101010101000001000011000100100010010001011110101001010111100011000110111001010000011011000010001010110100000001001010010001111111011000000111001111111101010011010111110011110000001110110111111010010101101011111101001001110100010001100101010010011010010100001011011110101111001101001001001000111000111001100101001011110111110111001100001010001011000010010000000001000101001001101101010101101000111111100011101001001111100000010011100000110011100110111000101001111101001111100011111011101000011101110111001111001010101011011100111011001110011111001100100101000010000001100010101101110011110011101111010110101101001110010111000001011111111001011111111011010101110100100101001110100111000110010000001111001000010011110100111111101111001011100101111111111111011000010110010101100000001110000110000011110100111000100000110011101111110001111101011001110010000011000011001000011000011000000000010101011111011100011011000000000100100011010001100001111011001101111010111101010111000001010110011010011111111000100100011010000001111110111111001000100100100010001100001010111001000101100110101110010100010000001110100001101010000010011111011011000111000111101111000101000111000000010011001101011010010001100011011111110110111101100100011101001101110100101011100010000111101010111011101111000101001111110101111000001000111011000100111011100111010011011110010010011111101010111001001100100000011010001010111011100110001000111101100101011011101100010110111010111000011010010011101000001000011010000011011110101110001111101101100010100111100110000001001000110011011000000001101000000110101110010111010101010010011010100000101001110110000000011001011001001010010000101111110000110010011011100011001001101010001010001001110111010110100011010010001000110110000011010100011111000000111100110010011110000001101100100110111011011111111001110110110011010101000101101110100010010011000111110010001111100001100110001010110100000010111100011011010001111010010011111111111111110110010110111111110011000010000110000110100001101001100000001010100111000110010111101111100001000000111000100110101000111110100000111001100010110100000011011001110001011010011101101100011011100101010101001011101101101110001101100011100000001001001101110101010000000010111100011111000001110101001110010011111010100010110101011001101100010110111100010011010101110110001111010101010011001000111010000110110000101011001001011011011011101011101010101001011011111111100111011100011000100010111010000011011011011011101010011010110010111001100111010110000110011001000110011100111001;
expected = 4496241;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);
#20;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd3;
noise_select = `BIG_N'b10111001001011100000110101101000011111011100000110010011000010010011010001011000101010110010100011010101001011000101111000100110100110000100110001110001110111100010000110101010100101111010010100110100101100101100010001011101011011110000110111011111111001100000101010010000101001000101100100101010000100010010011010011010110101111010001101000101001101010110101011011111011010000011001101010111110010011110001010010011110001110001011011101011111110000011001101110010010000010010011110100001010000010101011011101001000001100111000001100110001001110100100101001000000111110011100100000110101100001100000000001110101010000011001010101010000010111001110011110100100000110111111011011110000001111011111010010110100010001010110110001100001101010011011100000100001110110110010111100100011110010110011110000011111001011010101110101001010110110101000100110011011001001110100010010001011011111111110111000000000110100000011100100101010000010110111001000101000111111100001100101110100010011101000010000111100111100001000010001110111000111100110000000111011101110110011010111110011110110011001111110110000111000001000100000100011011101100011001001110110101110001011101000100001000101010110001011100001001110101001001001000101000000000001001000101100000101001111110111101001000111010011000000111011001100100101110011001111011101010001101101011100000010011101101100010101101110010111011011100001110100010111011001100011001111010111101101100010011110010001100010100110010000100111001011110001000001101110100110110001101111010111100011011011101101110101100100101000001110010010011011011111100111001110111001100100001001111000110110010101011001101001011100001110001100010000111101000110010101100000110110100100101011000000101111011101011001111011101011010100011010000101100000111111001010010100010011000011011100110110000110001000100001101011111101101100111011110111111110001111110110110111100010110000000111111111000000001100110011001110000010000000010110111000010101001100010100001011101111110000001110001001001001000011100101111011110100101101010100010000110010011001101100010001000101110010100111111001011000101001000101110110111101110000101110101110101000111011011001011101011001111000011000110100001011111100110101010010110111010100100111000000101100011111100110100011101010101110110000110001011101001111110100001100001100111101101011111000100101011111101101101101001101010110011010110110101100010111110010011100000011100100010100011010100010111100010011100000100011110011100011110111101001000101011010000101000111000001011100011110010010000101100110110001000011111001111100110100100111101111001011111001101100100111001100000001001110110011010101011011100101011000010101010100111010010101111101101001000001011100100001100100001010001011100010100111101000001111011011001101100000010101100110010100000110100111110101100001010010100100110101000000100011010010100111010101010111001100101100101001110011100000001101000100010101110001101011100010111000000101111110110101100110001010000100100111001101000100001000010000101111110000101101011110101111110110110101011101000110000000101000111000100110010101001001101001111000011000011011001110000101001011100011010100101111010101000100101100001100001100000101111001001110000000000100000100010100001101110000101100000011110110000111011110011001001101100100010110011001101100001000111001110111010000000110010110010101010010011000100110110010110001000000001011111010111111100110001000101111100101110100010010000101000101111001010101110011000111110010011001101110011011100110110100000111111011001000111111001100100101111001011000001110110010001001011011001111000101001000101111100010001011000001000111100011100011000010000011111001001000000010000111111011101010010100110001111101010101111101001011011110010111000101111010110001011000001101110011101110100010010100000101111100111111000100010101001110100100110101111001111001001111111111111001010100000110111110011000111011100101011100000000000111010111010010011001111100111110000110101101100101110100101100110110101101100010110001101000111000100001011110011101000000010010101001100101000001101111100101101011010100101111101110010000101101000010101000001011101101011111001001111101010010111000101011001011011101111001101011000000100011010100011110101110101000110011100100001101001011100101100001000100011100000001100010111100100011101001010001111100101000011100111111010111001010001011010001111101010100010000011111011010110111000011110100100000011111001000100001011111110011110111010001011100011011111010101101100000111011101110101011000000110001010010100100001011111010100000000001010001011100100011010101111100000001111110110010001010100011010101001000101001011000100101100011100010101000101011010000100011010001110010001110101111010001111111101001111110100101011011100000111010000110111111010010111001000000101111110000100111011010111011010110011011000011100011011100100111111010011110000001101011110111101110111000010101110101001100011100111101011111001011100111111100000110110101011001100111110000000010100100100100100000001101001001000110111010010101000100100100101110010100101100000111110111111001011000101110001000000101010110101000011110101000100010000010001100110010110010110110110101110001001111010110011100101100011011001011001111010111010010010010010001011010100001111011110100000011001110100010010101001100001111001111010010000011111101001000100000100100110100110010111011010110011111110001111100110011110001100100000011000110110101010011100011101111100110100011001110110101100111001000010110101000001010100111011101110101111010010011000110100110100110101101011101010000010111110000100010000110110010010101111101100110010000011011110001011101110100111001111011010011001100110100001111000001010010001010110111101010100000010010111111110011001111111110100011010101110010101000011010101101100111000100110100001001000011000100010101000010011000101001101110001000100101111011011100100100101010000111100000000010000110101011110111101111101111111001110100010010101110110011011110000000111011011010101011000000010111000110010101111110101010011111111010000010110100111110011110111000000100111111001111010001101010100111100100000001000100001000011100100100000010110001110010001101000000010110101010011111110001001110111010100111011010110101001010001000001001110111001111110011010001000000010100010101100011100111110110011111010001011111101110000100110110101100000111000110110110011011101010001101011011111111000010011011111110000110001010001111110001;
expected = 16009297;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);
#20;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd4;
noise_select = `BIG_N'b11010110111100010100001010101001011110110100101101011110100010010011111110111011010000110010000011010001111111110010100100111100000101000101011111111110011010100111010110110101101101110000000010011000100110101110101001011011101111101011000010100010111011101001010001011111010000000101001110111001111110001101110111011001111000110100010011011100100111100101101100101011101101011100111111001100100110010001000010010111111111010010011011001100111110011101101011110010101111110101111111110100010011111100110110101101011011100110000110110100100111101110001111111010110001111000000011001110001011100011000111010001110111111101110001001101110001111101011111101010110110011100101111000011001001000110001011111010101100010000010011110111011000000111010001101111010110101011111111011111000110111100000011101000010100110001001010000110100000011010101000111100110100100110001001100001011001101100000100011100111111110101010010010000111110011001110000000101000101010100011000101101010001011111100100101101011110101101000101011101011000101011101100011011011110000111001101001110000010111110010111010101111100011101101001110110011111001101000011111101110011110010010000111000011010011111110011001011000000111100011101101100001101001011101011011000000110010111011111100000110001110011101111110101001000101111100010101110001111000010000101010110111111010010110000110001110100101110111101001010010100101101101001010010011100011001011100101011000101001010100100011100001111100101000010011011010010100110100100001110010110011101100101101110111011000111111000001101011000010101101100011110111011010110101111010111100110010101111100110011001101111101100011010001111111101100111101100110101101010110011110100110001110011110010011101111011110010001110100110110110000010111110010100000001000100111001010110001100100001000000001010111011100101101110100010100100010000111110110101111101100011001001010100000010111001100000010100011101001001011100111001100001100101010100010111100110010001111111110101111101011111011001110010101101011110000000100000001010001110000100101111000000011011101001010110000100000011101000100110001000011110010011101111011101110111100000100010011110000001110111111110011111101101001111010110100010011110101110101100001010011110010101101011101101011100001101001100010011101000111111011001111010000010000110010000110100011010110000100111011011001010010011010110001101001110100011010000010110000111010100110011001111101100011000001001010000100001111011110000001111111001000000100000000010011011010110110110111000000110000000110011111001111111011000001010111100001011010000010010111100110011010000010101010111101111010011000010111101011000000010000110011001110101001110110100010100010101001000110100101000110100100110001010101111100100010000000001011101011000011110111010010110001001100001001101111000100001111010100101000000111011101110111111000001010100011111111001001010110101100111011100011111101100101011100110101110101111010111110001010110011110111000111011010000000001011111111111111100010110101100000111110011011010101000000101010100111100100000001010110100001111111000110101111010011011101100101010011001010001111110101010000111010100100110100000100101100011001100011000011011000110110001000000110110010101111101110110010101011001000100110011011110110110100001011010011101010001011000010110101111001111101110100010100011000100101110010101100101100101110110000001001001010110110101001000110001100111100010111010001011101010010010011001111000111100110101101010010000000100000111101111001001110110011111010010110010001010001100100100011000100011110011101010100110111001011100010111001001100111010101111011101101101101000011110111001000110111001011000111010010101111101111110001111000000100111001000010011111111111111110011101100010001101010101100001010100010001101010101001001010000011000111000010010110010110101110010101000101000010000111110100011000000111100111111010010100010110001110011111110100111101101100100110111000000001000000001111001111110011000001010110101101010001101110110000111111011110001101110011011111010100010010100111101010101001001111111100111110011111110010100001111011101000101101110010011101010100101100000001111010001100001111010000101111100111101110010000111010110100111001100001010000100000010001110011101000101100000010001111001110011001111100001010100001010111000101011111011100100001110111100000100001100100010110111100000010010100000100110111101011011100001111000010000100001011100001111001001011001101010001000001101110001111001101101011001100011101111110010101001110101000100001001100101001010000011100010110111011110000100110000100000011100111110010001011111001111000111010011001000100100111001000011111101011101000010000110010011001111001011111000110100110001100011100110001110010000000010110011111111010111111000011100100101100001101010100010010000101111101101100010111000101100110001110011000000011001111011111101001010001000100110110000100001101000011000100011000010000100100101011001100101010001101110100111010100111011011011111011111100100100110011010010011111010100010110001010011001011100000110010001100100000010111010010110001101000010001101011010000000001110001101111011000001010010101011000100110011101000001010110001011101010101010011011111010101110001010011011111001111011011100011001010010111111111011010000000001011100001011011111011010001001100111101010100100000010100001101011100000101111010101111110010010010101011001111101011011101011100101000101001001100110010001011000110000001111001010101110011001101010010011100100001101011101000001101001111010100010110110010110000011101010100010001100010000010011001001110000001110011010010000100010110010010110011001001011111111101111111001111011100011001111010000000010100000001110101010101001010111001101110000001100000110001100101111010010000101100011110011001011010101000010110100101011110000110010010101001010011100011110110100001000010010011111010000101001011110101010001001101110000001010100101111010001010011101000111011111010101010010100111101100010100100000101001110000011111100101010110101010011000000111010010100111011001100111100100001111011001000010111001010100101100100010111110010100011001010001011010000101101001110000001101001111001010010100110111011011111101001010101101110000110111100111000011001010110001010100101110011000001100011101101011000010010001111001011011010111001101101001111101101101010111110011011011001110100110001100101001011011000101000110101001001100111001011000111101100100100010101001011110001;
expected = 4589000;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);
#20;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd5;
noise_select = `BIG_N'b00010100010010001111111000101111101111100101110000100110111010111100101110100010100001101101000000010111011110100111111001011001100100010001011000100001001111000101111111110011011100111010101011000001100110010000110011010110100010000100111110111000100111001001011011111111001011011001111001100001010001111101110011001000100011010100110110101101000011011011101000010011010101101100111010110100111001000111000110000001000011110000010001111101101001111010110010110111100010000110000110001100011110010000010010110001011001100101001111100010101000001110011100011000001110000001001000100110011001111011101001000101111100000011111100010001111000110000101011100010110101100101100000101111110000110011011110001001100100111100111000111001011000110011110000101001011111001111101000111110101101101011011010110000010001000000010010100111000000101100001101010111011100101101001111001110001111110011110010001010011110001001111001010110011010111010101101100000010011000010000000011100100011000100010011100100101000010000000000110110001001110111110100001101001000111010010100101111010101000100011100100000111101111001111000010001011011010110101101110010101111101010100101101010110000001100111011010001001111001111101001001001000010010111111000011100100000010100110111110010110101111011011100010000001011010110010101000011011100000101000011100110110101010010110010000011110000111010001001101001101100010010000101100000011010101011100000001001011100111010001101100111111001000110001011001110000110010101110110011110111100101001110111101001110101000101100110011101100110110000101011001100010011100110001111000011101110101000001111101000100010000110111001101100000101100010011011110101101101010001110111010010001101100001000111110101000101100001111011111011111010000100101111010001010001001111100101000100001101100000111100000100101100101101100011011010110110101110100110000011101001001100101011110111111011011110110110001011011101111001111000000010111111110010111000010011001111110000011001100010101101111101001101111110111010010100111001010111010101000001110010111011010111000011001110101001000101011001000000100111100011001110010000000001111110000110000111010001000111001110100000000000010010001111011011011111110010001000100111010101110011101110110101011000010000100101100011010111111100100110111110010001010001000110111110100000011010011010111010011010111101110101010001000101010101001001000000000110100100101100100000111001001010100010011001111100111000011000001001011111101100000101011010011111101110100110000110110000111111011000001100001100010111110011001010110010101011111000001111001110001101101011011000101011111000010100110110110111011011100110110100011000101111010011011010111010001110110001010010010011000001010010111010100010110111001100111100101100111001001101101011010100101010110111011000100010011001000100110101101100000101111101011011000110111001100100001101010001110010100110001000100001010101000001001101101100110000100010110000000011101100101001111100010000001100000011010001001111111100101000100001001100010001000111000011010001011100110100111000011000100000101000101001111011001110100001110010001110101001110110011110000010110101101001101111100111100100100111110111110001011001111100011010100100010110000111000000001110101101000100111010000111111110100011110011110111011100111101001010110100000100001101101111100110111001010100001001000011101001011100011011001101010010010100010000101000111111101111111110111110100011001101010101010001110100010111000101010100010100001010111100001001011111011011101000111100000111101011101011011100000001010000000010100101000010010111000111110011101110010110110110001011100100000100011100100011100101101100011101010011011010101101011111100001000111010000101110001101100010011100000001111000010111010111001010010100100000100100101111100100111000110000100001000110100000101001010011101000100011101110010001000111111010000101100100011100011010000000001001110011111011100101000111000011011000011101101101000100110001100000000000000110111011000110100110011000011011111010010000110000100000001110110101001000101000000011000000010100010111000000001011101001010000011100101000110100010001111001000010110110111000000111011010111011010001000011100000100101101111011110011111110001110011000100110110010000100100111001011000011001010100000111010000010100111100100010010111000010001101101011110001000011101011000001011001100000010011100000101101111100001010111001100001000010110110001001000100001011011101010101101000101111101101110101101010100010011010011011111001010000111111011100000001101111101101000001101001100101010110000110101111100101101101111001101000101111110110110000001010111000010000111100001110001011110111000101110111000100001100111100100100000110110101011101011000101001100010100100011011001010111110111111110000110011000101010100001111111010001010010110100111011111011000011011010101000111100011101001001011001010010111101100011000001100110111100011110011001100000010110010001010110001100011101110111010110000010001000011111010101011101101001001010011100100001100101111111110011101110000101100100000001100101001101100111001000010110101001010110001010100100010000011110001101100101110001011111011111011010111111001001100100000010010100010000111100111101010100100111011111110101101110110000101101111101111010101011100110000111110100010100111101100111100110000111101001100010100010010100111111011001101001011011111111110111110010100111001111000001011011101111010010001101110011001110000010100110010000110011010010110111010100101111010000111001011011010011010111001110010110001000100111100011010101010111111101111110011000110000111101010110110001001000011010110000101010101111100010101011011000010110000011110001001110011100100111110001101011111000100010110110010001000011001010011001110000010000110110100010100100110100000000010110110110011111110110110110110000011011110011101011000001001001010011010101010001100010111011101010110101100000110011010000111010111000011110001100111010101001001110111010100000100001001100001110100101101001111100100110110111100110000110111100010010010110000011100111101110101110001001100101001101110010000000010101011001100100001111111010100100011111110011101011000100100100110110111100010001110111101110110110101101110010101011110001011101101100100011011001011101000011010010111001010100011011101110011001110011100001001010111001100011011111000001110001110011001010011111100111100001011111100001111010111110111010101000111110000010000111010001110001011101;
expected = 8023960;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);
#20;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd6;
noise_select = `BIG_N'b10110011011110000101010000110101000111010111011011101001001101110100100111001011011111110001111100010111110111011011101000111101111010011101000001101110010000010000101011110010111100000111011101011001011111101011100110100111111000011011000100010011010111011100100110001110001000001000011011010011000111011001011101010110110000100111000000101010001110110100000001101100110111011010100001001011110110111111101100011010011011101011110100010000111111101111111010100100100010100100010100011010110011110111001010001000011010000011111001001111111110010110100001011110010011010011011000010001000100010100111010101010110111011110000011001000101011000011010001101001000001110101110101001101010100001111000111110111111010000001001000101010010010011000101010011001000110101000100100111111100010110001110101010001011101010001100011000001111000000000110100000000001111111110110000010011011010000110010110101000110010010001011101001110000001100100011111000000110000110001101111010100001101001001110000111011110001110111100011001001000101111001011100010111000101001000101100110110011010111100110011000100011110100111000001001101100011011010010111110110101111100100101111011011001100011101100101001100000101000000010000001011001000100001110100000011010010101010111000101001101101100110111011011101111110010100111101110101001110001100100111100100001011111111000001101000101010011011101001001001000000110000101010001111101100010011111100011111111110111101111010011111111010110100111001110001000001101010000010011011010100100011101001001111011011011101011000111111100111011111111110100001010100110001011011111000101011111011101001000111100010010011010111011010000010001011010010011001101001001010101100011100011111000011101101100100011101111101111011011111000000000101100000111011100101111010000011010011011111011000011100011001111100001000111110111011110101000001001000101010001010100111110110001010100100101000011111110010000111110001100111111100001011011001101010011011001111101101000011001111100101111100010001011011101111101010000001111011000111011100100110111010111100100000110100100011110001010010010001100111110001111101110011110111001010101001111101001001001010000111010011001011010010011010101101000101100011001000101101101001111100010000001101000011111001110110101110000111111100111001001101001111100010100000011100011110010010111011000001010010011001100010001110100110010010000010011111011100111000010001101011011011001100100010000010001111111000011001000100101001100001001101110010001001000110101000010011000100001111111000011110111001011110111010110100010111101001000101010000010110010100110110111001111000010001100110110111011110110111101111100011111010000001110000100001100000010011100111001000100101101100110101010100110011010110111111111101010001001010010101011010101011010001101101011110110001111100010110110000110001110011000001001001101111011000101000101111100111000000000100011010001100011111011111010110100100000110111110000010011010011110111110000000111000110100001011000110110101111110011101111100111011101001001010111111101010000001000100000110111100001110110110001011011100011101110100001110011010100100010111000010100000100010010000111110101000010001110011100101010111000111011100000001100001101011100000100111000011111110110010100000111001100101101001011111010101100100101000000100010011001110010011001111111011011011010011011010000010011101110111001101010001101000111011001110101110101101010100101100100111001100100000100100100110111011001001100110000000100111101110010000001101111010110110111100001010110110011111011110011110010100000001010101000110011111000110010100010111100011100101101010010000011011111001001101111100100111100011111011000111011000110111101001001101001101101001011010001111100101101110001100100010111101000000010111001011001000011001100000001111001100110011010000001001000110011110110101000010001000001001011010000110010110001111110000101010001101111000100110010010100101110110111111100110100011010111011010101000110110001010110001010100011100111111011000111100001000100001010010001001101101100101101110010101100000000111001001111011000010001010001000001111010101111000100101010101100111001011000001010101011111011001110100000101101100001111011111110010011101111110101100100000001001110011101101111100100001111100010100110001100110010000101111000011000111001010001000110010011110001001010110100000110000000111001101101110110111000111111100000100110111101001111001111110001111111011001101111100111101101010101110101101001101101010011111011100101110011100001100010010011100100000110000000000100110001000111010101000110100000000000011000001101110000110100000110100010100111101010000111100110011101010011110000001100100011101011110111110101011011011110011100111010000110110100100000111111001001100111110111100111011011000110110010011000000001111010110000011011001000111010110011111110011001010110000000001001000001011010100001100000100001001111001011011101111001010001010001100000111001100001100111011010110010011000011001100000111101000111010011001110001111010100100011101011001100000011111010000100111011101111101001000001010010101001111011010101100001111100000011001010011101111111010001010100110100100101111111110011100011010101110001111000011101000011110000000001000100010111010100000000110010001010100101101111101001100010111110010110010100011111011111001001000000000111000100111100011011010001000001000100010011101010000001010100101111001110100101100011010101001010011110100011100011010010100111000101011100011100011011111000001101010110101100100101001101000110001001110101111101000001110000100110010010001011001100101110000100111000100010101010010100010011001101001000101001110000000101111110001100010010111110010000010110001111011001110000001011001000101111001101011000110111101011111010001101101011000111110010111100100010101000101001101110010110000011000111110111011111011011100010101001101001100011110101010100001000010001101000011000010111110110001000110100001111011111100101110010001010101111100110101101101100101110011000111001100100111111011101110000111100001010010101100011101001011100001001111101100001010010111001000110100010100110100100011111111101101100101000101101011110001000010010001000011110001001101100001011010010111101011101111010000000000111011100001100010001010001100111111001000000000110010000101011110001010001101101010111101000100001100011111011101011101110101111110110100010110101000000000011100100110101101110110110010101100101000001111010100110110100011001110011;
expected = 7680713;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);
#20;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd7;
noise_select = `BIG_N'b10001000100001000110110110000000101000111100010110010111101010000001000010111101111000000011000101000001010110100010011111110011011110100001011000100010111001101000100100000100110110011101110111010100010011101000001101010000011000111010000010001000010011010110111101000001011000001110010100100011110000010100000000011010001001011011100011000110001001110010011010000101010100011100000101111110101110110100101001110010100000011011011111110110111100101101010110010110000101011110101001011001101001101101000101110110110110011000101110000110000000000000101100010000100010101010010100011110001100110100010111110101100010110111100011101101000110100011000111110110111011010101011101100100101001000110100001111011010100110111011111110110101011101100010100001100101100010001110010101011101110101101111011111101001100000000010011011101001011101001000001111111111110101110100010100100011000011010011011000111000111010011100101110111010111111111100101000000001011111101100010011100010100010100010110010010101111100010100011011101010010110010010110011010001100001101000001101001101100111101111000111111110100100100011000101110110001001101111001010010101000110100000001001010000101001000010110010011111000001101000001110100011110100001100110000011101110111101000101011011010111011110101100011111110011110111101001000110110111000110110101101001010000011000011111110100011010000010100010101001011000110110000000110010110000101000100000011101010000100011010001001111001011001110100011010110011100100010001100110010010111000110010001000101001010101101001101000100100100011101011010110011110001110010011110011100110011111010011011010110000100100010001111110000000101101011000010011010100000111100110100111110011101111010100001010000011111001001010110011000100001110001111111010100001100001101110110110000101000100110101101100110101110100100111111110101011010111011110010111111001101100111110000101111000110101001011010000001100000101011011111110000000000111111011001110000101100011101000111101111110000010110010101111000111101100110101001011101101010110000001010101110110100111000010111111000100101100010001001001011001100011100011100110111011001101111111101101010101111101110101011011000011010110111010101011110011010101001011111101110110100101000010110000001010100011011101111011111100101111010110001100101010001001100110111101111010001001000001100111100111110000001101101100000011001111010111110000111011101011001100101000011101011011110010101001001001110111011000010100110010001000110010110111011110011100110111100111001101011111110010001000001111010001111001011110001000001011011001100010111111101110111010001001101010110001100111101011010110101111101101000000101100010010001001010100101111100111101101111111101001110101111000010011100000000100001011000100001101001111101110100111111010100110111110100011011011011100001101110001101001011010101110001000001001000011110110010110000110101011000000000111110010001011101111110010100001111010111110111111111011000011111110001110000010111010110000110111011011001001011100111011110111110101111111010101110110001001111100010110010010011011000001010011010001111001111111000011001000000100100100011001100011100110010011001111110000000000111011001010001001100111001101000010111110000110110001000110110000111011101100011000010011100000111001011011010010111000111110100011110011011111000000011000000011101110100101000001010100100100011110111101011111100010100100011110011010010010110101111101101010111001110011111100111110000001000010001011010001000111010011010001001111111100010101110100010000101000111011011111000010011101010001011100011001100011100001111110110010011010010101011010000100101011110011111100110101101101110101101001110000100001110111010111000110011111111111010111101100011100001110111001100010010110101000001101001111011011111110010010100011001010001010011011000101111000110001101000010100011000000010111110101000000100010011010011010111001000010100111010100111100000111010110110011100100001010100101011010010110100010101110011110101000111010101101100011010010110010001110100011010110100111111000100100110111101011011000000001011111011100100110011100011101111101101111011011100100100001100001101100010100110110000001110110101101110111011010000110001110011001001010011100110101001010100101001101110100011010101100000110010001100001001000000111110011001101011001010011000100111100001011001010010011110001001100110011111010101100010111010011101001111010111111100110111100000111111100101010010111100010011010001010100000000001111100000100001101000100000010110100101011001001001111000011110011001110110110110011100001101000011001001010000011000110010110000110001110110000111111100010001110010110110100000110001000010010010011101000000010111100111111000111000111110000101000000001101011011001010100001111101001100000111000100111010100101101001111000010110010000000000001101100001010011001011100100001001011001010001000111101001111111001100111111011010011100111000101010010101011101001111111000100100111011000101011011001001111111000001011110001111110100100110010000000111000100001010111010000100010100101110110110111010100011111100001011010000101000000101011010000010111001111110010110110000011000110110101000101101011111000000000011111001001100000011000010000000101100010100101100000101101010111001000100001001101111100111110010110001110111010011001011101000000110011110000111000001101111001100100001000110001110101100000000101011011110010110001100101100110001111101111101010101011011011110011100000101001010000100110100111100011000111001010100111011100011111111110001000100010100110101001111100000000100110011101001010110111111110100111011100111010000100010110001001001110111111110000110101010000101100010101101110100101011101100010011100111100110001110101101111100110100010000101010010010011101101001001011011101011101101100011011010001011110001010111000010101100000101100001100111111111001011101000010010110101111110010101100010001101001001010001100001011010111010010110010110110111011101011001110011010111111000010111010100111101111011101000101100111001010101000110100001011101100100111000111111010110101111001011101100111011111010001100111100001100110111101010111010011010100010110101000100000000101110000100010100001101011110110010101010011101101010000001101011011001100000111100001001100100111101100100111010011010110110110011110101001100011010010010000111101110111011010000000011011110010000100000111111110100011101100011001011011110010011100100111000011110011001001100110100001110100;
expected = 3754740;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);
#20;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd8;
noise_select = `BIG_N'b10011001001000100001101111000011010101111110101011010100111111001000001110110011111010110001101101110000010101010101100001101011110000000101101010101001100101100010010111110011010001010110001001001000010000101101000111111011101010110100101001000110011001100001100010100010100110100010100100001001111110101101001001001011001000011001001100110110101011101101111100110001000111100010000001000001101010100100011100000100011110001101010010111010101110111001100111110101111011001101110110000000111001100100100000010010001100110011100001001100101101100101011010010000110110010111010110111011110101000001010000000100000101100111011011000011101110100011001111111110101110110111001010001101111011011010111100100010100111000001001110011010111001101011011101110111101100001101101100001011011010000110010100110101100000001110011101011001111011101000100101101001101101111111001000101110110001100011000011011000010101010100011001100000110101110010100100001000100011110100000011111011110010101100101001011001001111001100100110001001111111000110100010100000111110110001001100000011101110110110100001100111011000000010100110001010010011010010101001101001100001001001011101001010100110110110001100101010011000100001100011100110110011001111100010000111110101010001000100110110101110000100101100110100101110110001000111101010110010101011101011100010101100101101011111100111101101111011110111110011010100001100011111110010110001010000010101000110001110000100100011111100001101000001011011101101101000110100010110011000000001111001110011111111111011011100000000010011010100011100011010001100000001101010101001110001111011000111101101110110100011101001010111000110101001011101111001101110000111100000110011111000000011011000011001011101000111100110100111100110011001010111011100100001000100100101010010110000111111011111000000001111001110110111010110100111111001011100110000001111010011101101110000011101100100011011110110011010010110111110111100011001101011010011000011000001111000001110001110010010011001101000011001101100100011101111111000100010101001011110101110101001001010010110011110000100100010100110000010100000000001110010010101100001000001101001110101000010100011101000111010101111111011111111010010101011100101100100101110101100100010010011011010011001111111001000011001010101001111010011010000010000100010011010010111011100110111101010101010111000011000111001010111010111000100111000000011010011001000110110000111111000000001110011000001101000111100111010000101010010111000100001011101000001110000010111001000010111000001111001011111111001100111110100100110001010011110000100010001011111011011010100111000011010111110000010111000111100001100000001011101100100101001110111000000111110001100101110111011110001101010101010100110001011010000111101000100001110111001000111001000101010111000000111010101110101010101100011010110001001001101011001010010001010001101101100011101001110011001011000001001011101110101000100011110100110001111011010100010111000000111010000100100100111101000101100101011010111110000110001110100010000100111101010001011001000010101010011000001100111011111101011101011111100010001100011011001100010011111010011000011110001000101110111000101101011110010011111111000100101110010001010110101100110100000101011010100001011100100100111010010111001010111110011111011110110010101001010101011110110010100110011010101110101110100111011101101100010111100000010111111111011111001110011000000000110100110111101011101010000001010001111000000010110101010000111000111011100001100000101011111000001100100100011101111111100000011010001110000001111100110010101000100101000100011010001000001000001101001110111010001011111011001001111100110110100011111000000110000011010110101111000000010001010000110100110110100011111110001111111011101010010101111101101111011001001011111111111010111101111101010100101100100111111101010101110101101011010111111100000101110101000011011111111011001001110101001111111110100100101011110001111110000111001011110100111101110001011010001010001100110110111100100101111011100000000010110110011111111011010100100110101111110101000001010010001101000011001100111111000110000111101000011100011111001110111100100101101011010001101001111110101010111110101100100001101011100100001001001101101010100000101100001111011110101100111001111111001101110001010101001011111110001011110001111110000011110111100011110001001100010101001111000111100011100000000010001101010101001001100110101101011011011111110110000010000110110000011110010011101110100100111001000011110110010101110011110011000100001000101001000110100100011100001101000100100010110011111101000110100100101111010011010010100100011101100001010111010111011011011111010101101101000000101011011111000001001011100011100101110100000000101000111010111000001111111001110011100100111110111001110000111110110000100011100010010101011111000001111001111001101001101010111011100111100101110011011100010010011101010000100011011010001010010111100001111011101110000111010010111000000110000010011111011000001110101110101001110011100001100110001100001011011101011111101011111011110100111001101101110100110100000111111000010110111001100101110101001011101010001001110100011111001100110110111101001011010001111001010110101001011110111110111001110011000000100111010011100101110011000000101011111010101010010101110101010100010001001001010011001011111111100000101011010100110100100000011011011000001111101010110000110100010110110010011100101110101100010001111110011110011000111100100001101011011001110011000010000100000001111001000010010101000111000100100101111010110101110100100010110100000110110100111100011000101001111101110100000011000011110101010101001001001110001010000000011111010001110011101100001010111001100010100111011111000011110011001101000001000101101101011000011111001100110010110101110011001000011011001001100100011100000000001010011111101010111100001001101000011110000100110011000000101101000000101011000011010101011111100100110000110110000000000011010001001110010010101111100000011110101111000100001100011000010000011001011101001001101110001000111011001111101011010010011110011011100001001010110101100011010010111011001110000001010110111010100100001110001110010110001001010011010101110001101010111001010101010101000111100100101000001100011011110111101011111111110001101011001100100111101111111111000001101100000111110100000010110001011001010101110100000000100011010001000101101110010010100011110100011110100101001100101111000000011101001010010100100001001010001000010001001111;
expected = 10671308;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);
#20;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd9;
noise_select = `BIG_N'b11110101001000011011010000010100000100000000010101101001111011110000000110011010011010011000111101100100011110100111110011011001011101101000110011011110011101101101010100101101110110010000010011011000011110101011101110011111100101110011000100110111110100000100101111001010110001110110001111111000111111011001100001000010101001110111111011000110001101000110110101011111010100000110111111010111100100011001010010111001000001101110010100100010100010111111011011000100111001100011001111100001010000010011100011001110000011111101111111101001010100000000101010010100101001111011101101100011110010111001001000000010011100010001101110101001000110000010101001100010000001111011110101110111101011010111111011010011011110110000000111001101101110000011100100010111110111001000101101011111111001001100000111000000111011001010001110100111010000000101100001100011011010101000101100011010000111111001001111000000001111000001000111000011001001010010010111111101110000010001101000011010000100001100101000000111101110001001110011110010111110010000001010110101100010000111001101101101010000111000111100001010001011100000101100101001011010011011110001110010000110011111101011101010110011010011110001110111110110000001110001010011111011110100101111110010000100011001100010010001001011101011100001001010001000010010100001000011111011100000011101111110001111110010011011101001011001100011100101011101100101110101011011001101100111101101010101100000010000001110010001010110101010111010100111101111011010011100100000001011010110001101011000011000011100110100001111000011101000100011010101111100101111001010011111001110100010010111001101001111011101100111000000011101001000011011100011010011001100111101100111001010110100110000010101111011100011010110001101001011110100000000101100001110110100110010110110110100000011011111100000110100011011011111001010100111111100011111101110011101010111101101110001000001101101111010110101111010000111101001110011110110011000110101010011111011000000101100011111011111111100000111010101000111010011000010011001100000100011011110001011100100111010101011001100011100101100111000100001101001110100111001100010010100010101001111101010001010111000001010000100010000100010010111100100111011100000110000101010100111110001001110010101011101011100001101100100101110110011110000010011000101110110110011001110000000011100011010011111011000111100011000100100111111011010110110011011011010000011111000100001010011010110011010101100101000110110111010100100010110110101010111101010011000001010101001010111101011101111001010001000010110010111101111010011010101101110010010010111000001011111001101110010101011111001110001001011010100010011100010000011110000010111111110011000111010111001000011000001010011101101111111000111001001011110101011100101101101010111010000110000000101111101101001010100000000010101110101000000000100100000000000100100101000010000000101000100110110011000010001001111001101000001110111000011100100111001000110111100011111010011111011110000001111101110000110010111010111000010111100000001000001101001100100101100000101111011010110101110001101001010001110010000110010111011110001010111010000100100111011110110111111001000110000111111110110011101010000000000111010000011000110011010010101001010011010101110100011100010000001111101111101110000010001101010111110111010000011010101100100001100110000001001101010000010010000011110110001010100011101001000010100000011100010101110010001111010101110100100000101001011110100100000111000110111111101111110001011100010001001011100111100001110111111101111010000101110000001111011001110111101100101101101000111100110101011011111101001100011101111111110000110001010100011000101111011100110101110101110011010001000010000000111110010000011000010000000101010001010100101100110110111111001111010100011101100111101100111111010010011110100010110100110111111101010011111001101010010111001100110000111101101110001110001011011001000001111101001110000100011010110110010000011000110100000000110001110001111111111100111000010010011011011011001111010110111001110001101110111011100011011000011100111111001000000111111001011010101011011110101010101111011001010011110011100100001111110001111101110010000100111101101000000100000011001100011101001110101110111111010100100001100110101010100110111111100101001100000100001110101101110100000011000001101110111001011101010101101110000011011111111101100111111100101010100011000110010010000101010010111110110011000110110000101001101111110000011000110010100101100010010101111110111111011010101110011111011000001100010101000101000100111011110000101000010011101101100101101010000101011000001111101001110110010110111001011011110001100000010111100000011100110001011010101001000000111111101100110001011111011001010001101111000110011110000011000010000110011011111011000001110100111000111001011001111000101000001100000001000101111001111010101001011000000010010101001111101011011001101001011001110011101011011111100011010011010111100110010001010000110100011010110110011010010001111011010101101101001111010001100001101011101111101101110011011001001110100110111101010100100111000110000101101010111001100001001100000001010110010010011011011111100101000010001100001001110001101100111110111000010000010101010001111001000001010001000101111111010001001110111110101000111011010100000110111011111010101001101001100111000000101100011111110101100110010001001011010001001100110011110101001110110110111010110110101010100001010010110101011001100001111101101000010000100000000001010111010100011001111011101101110011101110100111010010111000000011111111001111111001101001110110011011011001010000011100111001010111101000001001011111101001001000011100111101011100111110000111011000001110000110001100100010110011100001111010101010111111010110001111011100011011000010000011001001011111000011111000001111001111100001100110111100101011110100001000101110001101010000010010111111100110100001110101101001100001010100001110000000001010010010010110101001010101110001101000111000101110010100111001000111010111000011100101100011010110100011110011011010011010101101011101100100011110100111111010101001001111110100000101101001111011011000000010000101000010101101010010001001111110101111011010110100000100010001100101010001001001010100100110111010011101100010110101111111100011011011101111001101010100101001011110111001001010001110000111101101100111111001010001011010110110001110111101000101000101111100111000111000001100001100110100101001111101110111101011001001111101100111010111110100000110;
expected = 13974784;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);
#20;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd10;
noise_select = `BIG_N'b11111010000001101100000000111100011111100011110111111010111100011011010000000001010100110110001110111000100000101111001101111101101100100011000001011001100111111100111100001111110000000110111001101100000110000110111000100010011011100101110010111001011010010100000000111111001100111101001110010001010011110011101100110000101100001010011001100011000110000011100110100110000100001101111101101101101100011101111111110010101110101000100100100101110010101001001010011111111011001111000100001100111010110000000011010001111110010000001011111000001000010100010110100010110011010011000110100011111000001001010000110001100011000101100110110110010010111001111010001111100010011111010100101010100110011100001111000100101001010000001101010010011111111000000001111011001101000101101011100000110100010000101100101110001011100100011110011100011011001110101100001010000000001000000010110010011110100001010011110010100110111001000011010001110011110011011001101010011101110101111010000101110000000001111001111110110101000000111011000101011111110100101111100101010100101110100011010111110011101000111100111111011100000010011000100000010010001111011101011000110010100000010011000111110011111010000001110110001011001010010010011111110100111111110100001000110100111001001111100000100111000110010010010010010011101011101011010101111101100110000011100010001110100001100111011100011011100110111001110010011001111110101001110101110011100011100010100100010001111101101100111100110101010101001100101101011010001001100000001111101101110100101000001000100010001001000100100111101011101101101010100001111101100011100110101001010000001100111110000000100111111000010001000101111011001110010100100101111110111100011100010010000010001110101011110100111010010011111100001000111110100010110011001111110000101101010100001000000010010001010010000001011010011000101111010000110011100011110011000101011101111010101100101111101100101011111101100001111100011000110011000000111000100011111001000100000001110001101010011011010111100100011110111000011010011111100110100000111111101000010100001110100001111001111101000111010010011010110001000110100000010010110010010010100110000011100000000100100011011001110000011011010111001011001100011000011010000000010001001101011010010001011011001001110100011000001101110011111110101111001000000110000010001101100000011000111100001110001101010100011100101010011110001011101111101000100011001111001001011000001001011010100111011100100001010001111111010010110111010110000001010100101001101110010111110000010011001000000101101101100110100001110001011000001101011010110011011001110010010001001001011110100000010111000100101100110011011111000101010011111010110110001001010010101000001111001101000010101000101000100010101010110110100110010010010101011010000110101111010010011111101101111001111101000010100100100111010000011000100000001111011000011000000100111111111011110010001011010100010101011010111011110110001001001011001110000110001010001111011001010111110111100011110110011110011101100010110111001000001010100000100001000001101011001100001110000111011011011101001011010110000101000111101001001011011011000100010101111010000011011101110001001111101000101010111001101111010101100000101001000101110101000010111010001100110111111111110010001001100000111010010110100000010001001010100010100010011001000001011101110111101001000111101110010111001110110111010111001110111010001101110100111011000111101001001100100010101001110110011101111001100010100101010011010001010011111100101101001101001011010001111000001101101011001101001111010100100110010011010110001000111001011011110000101111110000010000001000000101001011010111111000110000100111100000100101110111110100111010010110010011011010110111100101011101100011110001101110100001110001111100000101110011110000101011111011111100110111101010000001011100001011100011111111111111100011010000001111111001010000110011000010111111011001000001000001100001010101101001101111010011101000111100111101001000100111101100101111100100011110110101111011000001101101111000100111101110110101100100101011001011010100011101111110100010010011000011110110101101011010011110100101011010100111110011011000111101001111011011101110111101110011100011111101110000110001001010011010111011010010000111100001000011001111011101110000011001100101111110111100110010100100110001010101101001101000110011001010111110001100110000110100111001000000100010100110100010000011100001101101011000010010011110100011101111001100001101001100001101111110011010101100111111110110110000010110001111010101000101111100110001001110100111110101110111100011110100010111010110000100100010110001000110011000001110010110010001101101110111010101100101110110111010011010111111000111010011100111110101001011101111000100011111001100110010101010101010100101010110101111001100111101110001011011110000010010111010100101101010011001000110111010100001000001011100000000011001000110011111001101001010010100110010000110010011010010001101011100110010010110011100011110000011001011011011100100101111110001110110110010110111010101111010001000111111011011101101001110001000110010000110000111110110101100000001111110100100100110000100010001110001100010010000010111011111000011111101100101001110101110000101110111000000110010101010100111010000010101101111010011010000010100111000011000100100000000100111011011010000001101100100101010010110100010001110111111000101100011010011011001100000100001111011010011101001101011011111011101000101110010101110101100001001001100001111011010010010000110111001100101110010010000010101100001101111011001110000000011001100101001001100100010110001011011111001110000010101111001001010100110001000000001011101111110111110101100101111100111100101110100001100000101110111110000001011010110001100011111100000000000001010010111010110110111100010101111101010101011010010111111110101100111001011011000111111000001010110101010011101001001111110000001011000111000001101100111101001100101010110001101110011101100100111011000110011010100010010110000110001010101110011111010101101100110010011011110100111010100101010011010110000010100000101100100010100001001111111101101000111110111111111011000111010101010100100010011001111101100110011011001110010100001010000101011001110100001101101001110110100111100101101110010001000011010111100000011011110010100010100100101101100101101111111111011101110100000001111010111000010001011001101111010101111010111101111000000110111100100111111111111001011011001100011111010011110011101100001111010110111110001011101100;
expected = 11462644;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);
#20;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd11;
noise_select = `BIG_N'b11111001010110111111101110000011100011000101101101100000100101000011011011011000001110110000100011001010000000101000001101101010001100100100001011000100010001101111001001110100100111110010011101111001001010100101011110001000010110000011100110111011011010011100000101001000110110101011100111000010011011101010001001010111010001000111000110111100100101101111110011000101101100010110010110100010111001010010001101001000100001001011111011011101010010000001001111101010101001111100010001000001001100011010000111001100110110010101000000100101111101111011101110111011110101110001011010010001001001101001111010110100100100000001100100100000011111111000110110111011001111101000001110100000011001110011111001111001110111001001100100010000010111011000011101010101101110111011111010101010111011010001110100101110101000110011101001011101011001010110101001101000100001100101111110101000010101001001110111010011000001101001111111000001110101000101001111110111101001011101111111100000011101100001000111000101011011110100110010001111101000011010010111100000101001011000110100001101101101011011000001000111100001000010000101000011011110110001110101111011000100001111111110111010011010010100101010001111010011101101110110001001001110001111101011100010111000011001101111000010111100110111100010001100110110100011001101101101010001010010001010101101101110110101110111111010111110111110011001101011111100100010100101101100010100000111011011011100101110001011001110111101010100011001001110101100011001001101011000010101110101101010100101011010011010001101110011111100011011010101111100100001010110010110101110001111011001110010001000010100101001111110010100101011010001001110000011010111000001011011101100010110000010111101011010100011101000011110010100100001010011110011000010010100001011100001110011010001011010111110011100001111001010010100100000110101011001110010011000001100011010110100011110011011110000001111000001101001010001111100100100111110110111101001111101001100001111011110001101011110101000111100011101100101110000101101011100111111011001101101000010010110000100000100000111001111001011101000100010010010101000111101011011110100010100010100100101010101010110011100110100000001010111000100100110101100111100110110101110100101000010100000010011111000110111011011100100010110101101101100101111001011110011010100100001000100101110101011110100010100000011101001100011001111100000100111000100000001100011100010010011011111001010011011011110110010001010111001011000101101000110000000111111110010010100011011100011011010101011110100101011100101001010000111111110111010010110101100100100001010000000011110001000100000000110111011000001001001110000101110011110110111000100001101100111111100011011101100101000110000010110001000100110101100010010111100110100111011111000001110110010010100110110111111001000101000111011100100000001101010100100011000000111001011101001111011110101010000010110010110011101001010010001001001011010010111110010010101110110110101100101000101001000100100110000001111101101111111000011101000011100110100101100010101011110000111110110111111010111110001011110010101000010110101001110000110010101011101010111010110001101000101110111110101011100001011101101010000001000001010010011010100110111010101111100011100001011011110000101001001110101000011110011010110000110001111111001000110010011001011100011100011000010111000101100101110010000011110011010010011100101011100000011010100011001000101010111000010001010110011101111011111000011011010001100001001001010000011110101010100101111100110110100010111100110010111001000011110011111011101011000010001010011011110100011010110001011000001001000010010000111001100101100111011110100001001110001101001100101011010110111011100000101001100110101011011010000001111000110110100111010101111010110111101100100000111000111111001001010011001111100100011010000001001100100000100100001110000000010000011111011010011110000110100100000101001011001011110011010100011110000000000101000011011101010010001101110011100011010001100010110001001111001110010010011111000011111111010001010011100010011100001111100100010000110011001101111010011100011000011110010000110100011100011010101001001000101101101111100110110010110101010100001100010000110011010011100011001110110101101011000110110101101011101001001001101110100011001001010000110101000101000100101111010000101011010101010111000100101110101101001101000111010101001001011001101001000110000011101111010100000110101110010000100001011011111111010111111111111101001100100111101101110001100011011011010101010001010001100000011000000100100000111101010011101010111111101101101101100111111101000101111110101100110001001101110000110111001100111000001111001011100010001111011101111011101101000001110111010100001111110010011111101111000111001111110001010010000111000010100111111110110111111111110111011001011001111111011111011100011001010101101101110111101110010100110100010010000001010110111010010011010001001100110000101100110001001100111111100011101111110001011010101110001010100001111110110000101111000111000010001100101100001100011111011011001011001010101110010110111111010100100001100010011000001001111100100011000000001001101100100100100100001101101001100010011101000000110000110111100101000110001110110000011000010010011000101010101110001011000111010110001010110111111011110011100111000001010000110101100100111011100000011111010111110101100111011000101101100011000101000001100100100110110100010000101001101100100111110011010000000011111111100011001011010110110001110110010001111000111001001111001110101001110101010101000010111010101000000010001001001101001001110010000101101100001100000001001101100111000110100011001110101001011110111100100011001111001010010010110110101110001000100110110001100010011110111111000100010001000010001111000111111010101100011111001110100111001010001001001100100101001101110011001000000010110110110100100100101001110000100000011000011010001101100101001010100100110100110110110001101001001011111000001011101011111110110100101011101101110001010101110001011110011011110110001001011111011100000010111110010110010100110101010101111001110000110101000110101001100101100000100101111000010011011011000001001110001101101111000010101110011110011010100010110111100001000011101101110111011111000000101101110101011100000111000111110001010111111111001111110011111110110000001000010110010100010101011101001101111011000001101111010111100001000111000111101001000110111010111110101110000000111001111001011010011101010101011010001010101001110101;
expected = 9096790;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);
#20;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd12;
noise_select = `BIG_N'b00101001000000110100000111000000101010101010001100011001111100111011000001111000000000000100001100100111111010100111100011011000010101101010000001001100011010000011101101101111010001011000010111001101110000011001101010000010010001110010000110010101110011101110011110000001101010010000010001110001010110000001101011101100111001011010110110001100100001111110000101010011001010111111100111100001010111100011100101010100010111111010100000001001111011100011010001000111001111101111110000110101110000011101001001010000000111011111101010101001100011110101110001111100100000111010010010000111010101000101111010101100101100111000100011010010100111100101100100111011110011101111100001110100000010000100010111001011110100111110110111010010011111011001010001101000111110100000110000111001111000101011110010101110110100001001101101011000001010011011110111001110000111001001101011011001111111001001001001101100010110110100111101110110101111001100101110111010101111110100100010010110110010110111100010001011111011010000110110101111011110110010100010110010111100001100101110000110011011000010011111111110011101011000010000111001001111111010010110100101001111100000000111111101011010100000101100000010010111000111000100001111001110010011111000101100001001111001110011011011110111100100101001100001010011100010101100100101110001100101111001000100011110010101110011011001101001101101111100110101111100000000100100111111000111001111001110010111101100011010100010101001110010101010000001010110010000110011111100100000001111011111100010010111111101101010100100011101100110111100001101100010001000000001011000111111001110100001010100010011001000100101100100101001010011010001011011111010111010110011110011001111011111111100101110001100111101000111010000110100011000110000010100001101110101010000011011100000011010101100011110100111111100000001101011000101000000010010101110101000011101011100010010010010100000101110001101100010110100111110111100100011101010010011001001011001000100100010011000011111011010111011101001111110100111001011010110111010100111100011001010000000111100111111110101001011100010111110110011010110001000000110101000001101011111111111101001000010001111000101000110011010010100010000001000100010111011011111101001010001100100100100100000001101010001000011011000001001110011101010101011111101101001111111001001010010101000101111011101001000001100010101101011001010111011001001001010100110010011111001001110010000000011101011011000000011001110001110001001010000100110001100010111010011000000010100010010010101110011000011100100110101001010111100010011100111011001000010101001000001010011100111010111001100010010001010100011101110011100101001110000010110111111010001101101010000111101101100000010111101011010010110110101101111100110010010101110110100011001001110000001000111001110100000110100111010110101101000000110000011101011100101100101101101110010111110011110110011100011110011010000100101101000110100100100110110010011010010100011000000001000100011000000100001111000001000010000110010100110111011100001111000001110111100100110011011001000110001101110011000101000001011000000101000000110101111010010011111111100111100010000111110001011101100010100011001000111110101000001010010010111000100010001010011000001000011111001001001011111011001110101010100110101101111111101110111101000010110000100101001100111110111100010110110111110100000101010101001001100000000101001011010011100010110000001101100101001000111110000001011011001001100100111111100001111100001011111111001100111110001000011111001010100101110100110110111110000111111110010001001101111101001010100101011101111111110101101000110000010101111110111110110101011010101010001100100100011111111010110111100111001001001001110011110010101100110000011100100011101011000011110110010110010001110000011010101001111010100110100111010100001001011101000000100101011010011110000011100101001100000110000011011000010011000001111111111111101100100011000110110111110000100111001101101011010100100001001011011000101110010111101000010101111010011000001000001111000011101000111000110001001110000011010010110100010010000111100110011011010111101111100011010001111001101100000000000011110100110000100010110001000100100001100101011010010111001011010001101110011001100010101100010001000001001010011101101111111111000101101010101101111110101100011010010101110100011010110001101101010001100011101011101001001111001011000000000110001010010101011010101111010011111101000001101110111111010000000111000001010101011011101010000000000011111110100111100101111011100011010111100101110101000101101010001011001111000111000110111011001110101011101011001010010110101100111110101001011111111001100011110001000101101011011101000110010110101110011011110101101100101011100101011110000110010110101001111101110010011011101111001010000001000110111100000110110100100001001111100111001010101000011010010100111111011000000101010100011110000000111101101110010100110001111000111001001011011100010001010010101111111101111001011101000101011011100001010100000000110100000001010100101001110010010000110101010110010110100000110101011111100111001100110000011101111110000001111010011000011101101001010011111001001011100110001100011000011001100100100100011110011000001001110010011011001101000100010100101010011001010000010000000110111111111001011001001111000110111010001010011110011010001110011100001010011101101011101001000100011001100000000101000001001000100000010111011110010010010010011000011110011010110000111000100000111011110000011110101010100000100100011101111110100010000000001001101000000110100110100011010010001111111001100010101101101110011000000111111010101110111001000100110011111000000100000011111011111111011101000011100100010101001000000101100000111010010100110100100011001100001110001010100001010100011000101111000000010011000010000010101011101101111111011010010100000100010001000001111110100001111011100010110100110001001000100101001000110101010111101100110111110100010101110001000010111101100011100000011000101101110110000111110101010010101111011011001100111010000100110110110110101100101100110101000010100100011010011010111001010000101111101111101011111100100011010001000001111011111101010010011000101101000100000111001010110110101000010111001101011001000100001011000000010101101011100101000000100001010100000010010000000101101110101111110001100000101010000111001001101111010000010111000010000001111100101011111011000101011100100110111010010110101101000110111001101100111111111001110011000111110011000000001001;
expected = 8739487;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);
#20;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd13;
noise_select = `BIG_N'b00001001100000110000001010101010010000110101010101110100111111101110111010000000101000000110100110100001011000010100011111001011000101000100000011011000011101011010111010011110001000010001000110100000110010111000100000110100101101001010010000010110000101001100010100000000111101000011011100011100001000011100111011100000001101101010110011111101001010111010001111001000110100101000101000100000010011010101010111001011111111011101000001011010011100010010101110001010001101001000001001101110010111001100011010110001111101000111011001010011000100011011101010010101111011011010101001100000010011100110000010010111110100111100001001101010110101111011010100000111011101010010001110010101001110100011001000011000100111000110101000000001000000000011110011000100010100001101101011111111110001111101111011010110000011011110110110100010010100100010100101011001110011111100100110011001000110000101010001000100100010111001100111001000110110100011010111010111110101010100000111011101111011011010111110000100100000111100101101100101111001000111100000110100111011111001000100010000100101000110001101100001011111001001110101001010011101100101101101000010000000100100101011110011110011100000001100101101111100000000100001001011100001110011010100011110111000110000010011110001101100100101011000001010101111101111101000110011110110110101111101011111001100001000111111100101011111001101001000000100101011110110110100110000111000010100001001000010000101001010100100100111101110100001110110000110011001011010110101001110101110111110011001110000011110111011001011010101100000111110011000001101010000010101011111010001011100011010000101000110000110100000100110101100011100101101101100101001110111001111011111111101111100001010110011010010010110100111111111000001100001001110011111000100110011010010010001111011010000101001111101110011011111011100001001110111110100101100110110000101101110010110100101110011001010111111010000000100100001101000111001100000011111000101100011111110010100101000101100110010000101001101011001000010011101110001010010111010100011101000101001011100000110000111110001000000100111010111101100010011000111000100100100110111110011011011010010110000011011011111110000010101101010111010010000110111101100101101110001001101111100001100101111001111100000010000110001011011111001010001111110110101010100111110100110010100110001000000100100010101111001111111011000110100001110100101000001100111011110001110101011001010011111111100011000011100001001000100010001001010100001101101101110001111010101011101000000101110100111011001001110101110100100101111001010011001000110011110100100011110110011010000011001011111100000110110010101111010011110101111000111110100100011111001000100001111010101011011000001001100010111110000101010010110011010100111101111111110110001010100110101111011111110001011111010001110010111011010010000101100011000010100010110001000110111100111011010010011010111010000001011010101011110000100010110100001010110000111000100000100111011001000111100001000100010111010001011011111110101011010111000000010001011101110100100111111001100011011110110111111001010011111011001110111100100111000011100011001010100000101111000110011010100100001100001111001000101010101110000011011110100000001011101100100000110100101100010101010111100100010010111000111010010110000010110010010011111000010001100001001011111100011100100110000010011010100101111110001000100011000000101101010010110001001101101010101011111000100101110111011100110011000001111110111100010000100110110100000111011010101001011011100110110101000011101001110000010100100101011110111010001000001000101110010100111011001001111111000001011010010100011110110011100000110111000011111001111001000111110111101000000001110111010010110011001101011001110001111001001101011000000111011001110110000010101101001011101111000101111101101000001111011010010001001101011011110111000001110010101110001111001011010000111101001001111111010011101101100110011101010111101111110101100000001100110001100010110110111001010010011011110001011101011100100110011101000111011011010000101100000011101000111010111011111000010000011000101111110000100110101010011000100110100000010101100001100010101100000010100101010010011000001000111101110011010100010101010110110000101110000001110100001101011001101101000110010011110110010100001100111000100010010010000000001100110101011010111011010111101101111001011010111110000111000000111001100100111011000101001101001111010011111000110110000010101011100111001100000100001010000111110010110110011110111011100010011100010001110110001011110101100001110010010111111100100001001101110001100000101010010100010110011011100011101011011010101011101100100110100001110001111101011100000111011000111100101001001101101100000010000100100110110100100110111010001101101111100001001000011100110010100000101110100011000010101111110111101100101111001010111001000001111101100010011010111100010110000110111000010000110110111010011110110000101111100100010110011000110011000010000111110101000101101101001111011101110111011011010011001010110110110100111100000101111001100010000111001000100011001111110001101001000011101111001010010111100000000111011010011000000111001110010001001011000000011000000010101000011111101011000101101011001110101101011000011011011101101100110011011000100100001111010110001010010100110111110000000100111001001110001010001010110000010111000010010100000100000101010010110000111011101000110001100100001101011101001100100001010111000111000001101001111001100001010000110101110100010101111000001010011000011111000011000000101011100110001101001000101101111000101111001111011110010110011011110110110110110011111101110011100001111000000001000011101001101101011001100010010001000111110100011001110110000000100010101000101100010000110101010000000111011110011110000110111000110101111011111110111101011111101010000000011111110111001001011011100001110010010001011001010110101010101000000101011001000110001011001010100001001101011001000011001110111111001001011001011111100000110001010010110111111001110110010110100101000000111011101000010000111100010101000011011001110100010100111110011010111111100111001000010101111101000011000111101101011100010101100100010110110100110111101100100111000011110010010010100100011110011010001111100110001011001100110011000001000000001110001101001001001010000010100000110100110111011000111101011111010000010100100101001010000010110100001011010100110101010101000110111000011000100110010000001101100101000010010110111100110001100010001000000010110000;
expected = 14496443;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);
#20;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd14;
noise_select = `BIG_N'b10000110000100100101100110011010000111111010010111001000111110010100000011001101110111010001101010011000101101000101110000100111010010110101101100110110011100100000111000101110101110100001111011100000001010101101100100010111011011101010100101000010100010110111001100000001000100001010100111110101010000011101110111111100110110011101010100001011110010111110010001011000101100000011100101011111001010110101100100111110011011001010001001001000001100101101111111111111100100101000110100100100110000000000001110111010101111110100001111000111111111101000010111110010100100010010011011000100100100110110011111010011011110101101101000110010000110000111111100011110100111100100101000100111011000000101001101101111100100010101001110100010110010101101001100101110001000101100010001100011000011101001000011010111101111111011001000001100111010000100111001110000111001101101110100000111000100101100100010010110000011001011110011011101111010000011110001011011100010000000101100001010111010001000111111101000011100111001110110000101110001001001000011011100000100010010000111010110100101101001000011011010000000101111101110001010101000000110100101010001100110111011111101011101111000111111000110111000001101000000010111011010000110011001100001010001011001010110011100111010100001111110110000000000110100011111101100101000100010101011100100011110000011010110110010011110001101001000001100011111100101110011001000101001010111110000000110010010001100110011001101101011100010101000111100101010111001111110011111011010101011111011110111100000110101001111101100111011010100010001011011100001000110100010001001001101110000001000101100010100011000011011101100101100111010001101011000001100011111010111111010010011011001100100101011000011000111000011001001101111001001011100111000011111011110111010000101011011101111110000110010110010111111100100110000111100011000101110000000101100011010001101010101110011101101100111001000001011110000101001001011010101100010110110011010100000011111001101011011000100010010111000111001100000111101111101110011100110011110111001010100011101010100000100101011011010000000111111101111101001001000011011010011110101000011110011111010010111111011101110110101111000110000000011110100011100001101100001100000110101000001101100010111000011100001000001011111111110000101111010100011111111010100000110010111000011110110111110011101110111000100011101011100010010001010000011100110011110001001000010001000111100101001100001000111001101111111011011110001010101100111001110010111110011010010100001101011010100101001110011011100100101110111000011000000110010010011000100100110111000111001110111101100111110001001101001011101010010100011011000100101100111011110111001001111001110011010011001001111101110000101000001011110100010011001011001010000000110101101000000101000101111001100110001110000011101100111110001011010001000010010100000110000101110011000011011101001001100100000001111010100010011110101111100011000011111011011111110011010000110111001100100011000011101100011110101001000001010111001111011100110111000111111010011010101100011001101010010010101010111000010111001111000110100100110101101100011010011101000010011010111101110101001101001100001011011001110001110000110100011101100101100001010110111100010000001111001011110010110101010100100011000001010001110100000010010100001010000110000011111110010000111101100101110100101100011001101101000010000001111001001101100101011000000001100111001111010101111101000110101101000000100000111001011011011100100001110110011000101100000001111001111010111111110000011010110101011100000100111011000011000100101111110100100010011011110111011001111010101101011011010001011010111001110101010010010100010100000111111010101111001111101110010010011110011111010011001010001000000010101110111010000010001000100111110011011000111110100101101111001001111010110101111100100100100100101001000001011001110110011001110011001100010011100011101001010001110111101101000111100101100100010110011101101101010110110001001111110010110010110111001111100101110010111010111100111111110110101101110011110100011001000100000100001111111101111110111011010001000111101010100101110101010000010011000110100101101010010011111011011000000101000110100010101001100000101010011000101111011100111101001111101101010011011010000100010100110001110011001111100011111011111100011001100001011011010000110011100000110010001101001000111011111011110000001000101001001110011111100010001000100000000100111100100111010010101011101101101111110000110111110011111101010110010011110010010111010000001001101010101111101011000011100001100000101100101101011110100100101111111010111101010100001100010010001110000110010111111001110100000001011011001000100000010110100110111011011111011111001011001011010111001100100000110010110000010111101000110010001100000000100000011110000001001000100001011010100000001111001101000111010101000111110010101110101001010010010010100100100001100111110100110001000000110001000101110110000011111001010001110010110011011000100101010110001011111010010110000100011001111010100011101111111101100101001110000101101011110101100100001111011101101111110001101010111010100000001001110100110011010110101001110001010011001001110010001110101101011000000110110000010101010110110101111100100111000000011100111000110110001010000000101110101111001101110011000010110000111101011011000110101110100111101001010000100100010010000110011010000101111101101101111111001110100101001100111111110011101011101101011000111100110110011110011101101000000110111011011011100111010110010010000001100011010101100100100111001111110110111010100000000010111111011001111101100001101001101001100011110011000100110110011010010000000001001011110111110111011011010111110101001011101100110111011000111010100101110100001001000100111101011110101100100100110100111011110000100011001101011100111101111110011001001101000100011110001001101111100101011001011000001100000000001000111111011000010100110011001110110010111001101000001110000000000110000011111011110011000111100111010100100100100111101110000111101111000000010010001111111111110111010111010111010101101111001011010000011000101000001000000110101011111000010000011100010011110010001010110010100000100011110111000001111100010101011000001101010000101000110111001011001101001001000001011100110101111100101111010111101000100001111011001110100001000010000000101000110100010101011001111110000010001011111101101111111100010111011001100000100110110101111111001011101101111101111001110001011001000101011011101110011111;
expected = 13448832;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);
#20;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd15;
noise_select = `BIG_N'b01101101010011110010001001001000100010010101011101110110110000110110100111100011010000011101001111110111111011111100101000101001111010110001011111001001011010000111100001111000011001011010110011010011110010100001101100000011100010110100100010110011111101010010001110110100011001010011101000010011110111110101111010011001100000101111010110010001011111000001110101001000011000111111000011110000011011110110010111011011001111111111000101111111010110100110001010110011010011010000100001100111111000000001100110110100110101001101111010111101111000110111110001000110100111100011101111011001001011100100100100111001001000110001001110000111001100010100011101100011110010100000000011110101010010010000010101010000011101010000011000000100000111001011010000100111111101111101101010100111000000101000011111111110110011011001111010100110100001010011010001010000111110011010000101001100101111010010011101110010101100001011101001000000001101000011100000010101010010001011110111010110011111110111001111000101011011111000011010101000101000101001000000010011111111101010111011101001110100001011010001010010011100011001001000000111000010010011100011110111011111000100110010011000000010110110000011110101000111111010100110111011100110111111100010001110000011011010111001010011010000000010011011110110110110001111100000110101001101100100110001000011100110010000101000011101110000101100000001001111010110011110101010010110000100000100100110001001111001111100000011001110111001000110011000001111100011000101011010000001000001000001001100001001011001100101010000010001110001011111011011011000000101110011010100011100111111101111000110011001001011000000111100100010010101100001011101010010101100111000110111010001001000110010011011000100110011000000100100011001100111101111110111101110010010100101110000100101100011101000100111000001100001000001101001100101111110111111110101010101001011111000100001110001100010000100011101111110011001011001011111001101001000010001110011000100100101101000011011011000010110101111010011100010100010101110001111101001111011011000111110000111111100101110010001101101111101001110000000000110001011110000011010011101001111010100111001000101101010101010100011000111111000111101110101100101001100111000110001111101000000111100101011011010010110000001101111010100011101100010110000010000110100111101111100100100010010111110000101000010000000110101110010011100100001010001100110010011010100101101111000010110111001010010001100110111100010001111110011010001010001000110001100110100001101000000001110101110110000011110100010010010010111100110010000001000110011001111110001110010011110110100001110011100101010110000001110110001110100111000101000000110010100110111011001100110000010100111111001111010001011100101100111011110001001100010001010010110011001010001111010110000011100010010010001011010000100100000011001000111111010111100110100111011110100111101000001011000001101001011010001010011111101101001010001001111000001001000100111001011010001011100000111101100101010000011010100011100101110011111010001110101001101110100111011111110100100000011011100100100110100101110100101100001111100000000010000001011000000000001000101010010001000111100011101101011011111010100110001111001000110101100111111101001111111110001111101001001110001001101110111100110111111101011001100110001111011011111110101001111000000110000011101011000011000010111010111001100111100010110100110111110010100000011110110011010100101010010010010110111011110000011100100011101110111001010101111000010101010110001000110000101010110011111100011011101011111100001011010111001001111001000010110011011110011110011001011001001010110010110000100000010000111100110000110100100010100101101010110001010110010010100111101001011000100110100010010111011100011011101111001000001011100100101001101010110111100111101000111101010001110001110000110101010010111100101011100101110001010100100011001110011001101101100101101111110100111110001101110001110100010011100100000101010111000001110010111010011001111111110101110011011001100001010000000001010100001111011100110011100111001101010100110000000100000100001110001110100111010000100000101101011000011010010100101001000111011011001111001100101110000010010011000110111110000110000001101100100011100111010100110010001100000001110111111001111100000000111100000011010011100010111010101000011110100110111000110010110110111100011010110110010000110111101111111011010111011001000110100100000010100101001011101110101111111000110100001011110100000111010100111101001111011001010000111011111011011000000110110010110101100111111010000001110011111010111101001100010110101110100111100011000001101001110001100101010111011111001111110100110110010010010011000010100001100101011000110000000100010110101001101001110011000101000001001000100100110011001010110101100010100111100111110001111100101011011101100111010010111101001110111000101111001100001100101101100111011100010000110001000110000110101011110001010010011111110100111001011010100100010111110000010101001110010111000100000111011101110010000011001001111110100010010100111000100100111110010100010010001111100110101010000111000110010001001100010011101001010100111010101111111011001100000000101001110101001000110001010000011100110000100011111101011001011100010011101101001101001100111111010110110101001011100101100010110001011001001100100010110111111011010100100110010101000101101111100100011011000000001100010001101001000000001100101110000101010100000110001011010110000111111110111111101011001001110111011000011001001111001101100011010100011110001011011000101111110111001111010110110000000110111000100101111101111010100000101101001000101100010010010011100111011001100111111101101010101110000110000100101010111111000011000111111010111111100110010011100111001011010100111100000100111100010001011010101000100100011001011000001101000100111010110001100010000101001001110110100100101100010100011111100000011011000011001010101011110011110101001001010001110001001010111111111110000001001001100101010000110001000010110000011010000001100111110110001001000111100001010001100110100011010011000100010101101100000110000101010010111010100011000110011101110111111010101111110111100100010011111111001000001101110111011101011011101100001010111001100001011100010110110001010011111101101000111100010100010011110101111000101100001101000100011101100100001101100111000010111110010100001000100001101010111010100010011010101011011010011110101000101000000111110011000010000110110001100010011011101110010001000111001010101101;
expected = 8893088;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);
#20;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd16;
noise_select = `BIG_N'b10110101010001110010100111111001101101010000010111001011011000101110110100101001001111010001010111101001011101000101000011001000000001111000000010100110111011011101100010111000111000000000110110110111110001011011101111100011100010000100111011100100100010111000111001010011010101101011101011010111110010000101110010000101101010001011110010101010100100101010100111011111011010110111111011101001110011100100011110111000101011011001100000000100100110011110000100011000110100101100010110011101001100101011110110010111011000010110111001010010000011001001010111001010010001110010000100110001111110110011011110001111001000000011011001000100000100101110001001000011110011011101101101101110110110011000011101001010110011001010100101111110110011111111110000001010000101000001011101100100010000100010011111101110111011011111001111110001110100010001111000110000101011110111001001010001000010111001111111110111011000000001111001000111011011000101111011001110001101100101000010000010100101101000011111101000001000000000001110110111001001101011010101010111101110110000100111100110100101110111111001110001000001101011111111010001100010111000100110100101001100101011010001100001010100000111000010010010101100101111000001000001001110011111011010010000010011001000101110011100001111011010101011010011110110010000011000100001101101011111110101110101001100110011001111111100101100101000100001100100011110010010100010110000101001100001110010010001110010111100010000011011010111101101101010011111011111001100101011100001101011011100110000101110110000001110100100110100001110000000111111010000100000101111011100110011000010100101001010001101110010010101011001100111100001100100001101110011100101110100001100001011001001000000001110100110100111110100111011010100000000111011110100101000110010111111111011101101001000010111110101000111011101111101011111011001111011100100011101110011111000111110111000101111000010001010000101100001110111110000010100100010000000011111100010101001000010111101111100100011111010111101010111100100100010110011100101010000111100001001101101101000000110110111011011001101000001101101100000010010011101010101010000010111011000110010011101011000000001000010110101101001010100111011000100000101001101100011101101100111000100001111001001010111010110000010001111000001010101101001010011010101111001010111110001010110111000101100101111111110100001001101001010111100101011100000000100101100100000010000001100101101001001011111010100110101001100100001100011011101001111111111110011110100110011101010010001111110001100000000011001111011000011100011000011000000101010111010110101010101110011100101110010100100011110110101100100001000000110011000001011110111111001110000001011100011000110101110111100011000101111011111101010100001001010111000100011111000101001110111000001111010110010011011000011010110010000010101101011000100101000010010100101001111011000101100010011100000010110111011000000111010110100000011101011001011001110000110110100001000110001110011101000000101010011101101011001010110101110011111010010100000000111011111010110111001001100000111111101101101010011000101000011100001110101100100001010101111001011011100110111100110101011011011000101110000111100101110110000100001110101010111101011100001000001100011011010011001001100011100111110100000110100110100010000010110001111110100110110111110101110110101000011111000011011111100100011001011110111110001110110011110111010100011101010111100110000100011101010100111011101010110100100111001011001011111111000101001111011001000001011011010000011001001010000001011110010100111000001000110111001010111101110000110100010101000011011101100001001111100100111101011101101010100101111111001010110110000100010110010000010010110010001110010111111111100110010111111111010010010101100110011010100011110101111010010000010001110011101000100100101100011110001001111101101100011111110001101010011110001101001101110000000000111010100101111101100000101011110100011110111001101000000010001011110110100100001011011010111000000101101011111000100001111110110010111101110100011111001111011100001011111011100110011001101111000011001101100111001110100110100110111101101100001100100111001100100111110000001010011010011101011111001011100011111100010110010000111011100000110111000000000000110011100011100001101101110000111101011000001011010011001001010111111011100011111010000010010100111111010010110100100111111001111001011111000110101000111100100101111011010011010010001100011011010110101110100010010101100011010010011100000111010110000010001001000000101010011001011011001110111011010011010111110100101000011001111111100010110100100010000000111100011011101110101111110000001110101001111000000011100110011001101111110110001001010010111001100011101101000000010011000011111000010100111001001101010111010001010101111100011011100101010011101010001111110111010000010100110100110100011011011111001000110001000100111000001111001100001000101010101110010111011111001111110100110100101001111000011000001110010010110000000110101000011111001111101111011010011101010001101000000001110100011001101001110101111101111111011111010000000100010101010101011011101001010100011110111000111101100001010010010000101010110110110000011010101101000100000110111000100101000011101110001000111110001101100001011101010001001111001111101011110111001011011111000000111000110001011110001100101000001100011110100011111101011100010001111010100011000110001101111010000000111000010001111000011000100000010011001010011101110010000110011101011010011001010001010000101100101010111011010111111010001101111011011000010101111101011100101101111101110101111010101000011000110010111111011001101100010100110011110011001110101111010000101000101101010010101010011100110001101101000101100101010100100010000101011111010010011101101000110010111011010001101010010110011110010101000101010001100110010011011101101011011001111110000111111011101000010111000111111100101110011100101111111010010000010011001111111000100000010000110110001111101011000011000000010010010101100001000101000100111111111001101110010000011000000111001101000010001110001101010001100011110100000011001011001010011010110010000110101011010001111000000000010101100010101100101011011010101000110011011111110001010100111100111100100111111011010101101101100100011000101000010100110000100101101000011101011110011100001101010110100011111000100010010110010101111101001100101011100011111101010010000000111011001010100100000010000100010101100010011010110010011011111110011001110101111101010000001000;
expected = 5941701;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);
#20;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd17;
noise_select = `BIG_N'b00011011111000101110110101111000000010010001001001011001111000000101000001010110111110101111001101001010100100011010111001001110111111100111011100001000101000100010100011111101100001101111001001010001000010110011011101100001011101111000000111000101101010001000000011001010001100010111111001101001100101110110111001011010111100000010010101010001010010100110001010000111000011111011100000100010011001001111111101101100000010111011101000010101110111000001100100101001110101110001001100100010010110100001110100001101111111000111100011000101011111000100101100100001100111111011001010101011100111111100000100010100100010000000011111010001110001001010101010111110000010110100000110011011011111001011101011100011100010001111011111111000010000011011101011011101111010011100100010101110110001110100100001001000000010100100010010000001110000001001111100111110100011001101001111010111101101011100110111110011001111110010011110111000011001101110001111001111011100011100100111011010011100110010110111011101110010111011000011011011000010111000001101010001010010111101111010011000010000111010110000011110011100001000100101111001101011111011110101010010001001011001110100110000000000010000110010001011011010110111001010101000011111110010011001000101100111100001011110111101111000110111001010001011011001001001000010110000001011100110110110000000011010110010110100111100111011000001010110100110111111010111001111011011101111111011101011101111010001011010110111011000110101101101101101001010100110010100101111100100110001111110000001000111111011010101101100000111001000000111101011101100001111101101101101011101110000110110000000000100100001011000011101000100010001110010011010110000101001000011010111010010101100010111011000000010001110101111110010110011000011101101001011011010011000010000110111100011000011001111001010001001000000000011001000101101111001001001110010111101001000110110111001011101110100110011011000001010000110101101011111010100111111111011010001111110010011011101100000001011011011111111011010010000100111110100010101010010110011010101111100101111111010111001101101100001101111000001111110010111101000111011011100110110000011111000000111001101101100101100001001010110101100010110110111011011101011010101111010001110011011101010001110011101111001011001110000010001000100000001111000111001000001000111110101010011111001110110010010100001100001111101010001110000110100011111100101001101101101100001000101011110011100111100011011000010011101111101001100011101101111110110101101001000010110111000110110010100000100001110011010110000100001100011011001110000011111110000001100001011011110100010111100000011100111110101010011100000100111011010001001100100110010101010011101101001010000110000000111101011100110110010011011111101111110000110000110110101100001101101001010001111111000101111111011111000000100101010100010110010000011011000100001100110100111000111110110000001110100111101101000100110001000010010111101000001100010001100001011011101011000110001100010001111111110111000110011110111111111000011100101111111000101000111100110111001000101100000110101100111001101001000111110110011001011100011000010100010100010010111100111100011110110111001010110011010001001000100110010100111001001101011000011100110110011100101100000000110100001100100011000101011110111000001011000111010111000000110010000000000000100111101110000100000010011110101011001110110000101101100000010010001110011100000111110000111000000010101010101010010101110001101000101111111111111111000101010111001011011011000100101001010100010111001111100000110011110010110000100010010100010011111110110101101111100010110101000001001001010011000110010000110101111110110010100111110011110001110010101101010000000000010100010101101000100010110100001100011000001011000011011000101011101100100000011100000110111110111001000110010100001111011010100100001111011011010001111001101011000111001010101110001100111100000011001010001100101100111011010111001101011101111101000010000001110000101100010100001010111010000101110111111011110110001011101110110001000110010011111000010110101100111010101000001011010010011101010100110111000010001101110111001111101010111011000101010000000100100110011010011000010111110010000011001011100011111110001101110111111100100101110100110101110110010000110101111000000111011100001111001010001100111000100011100010100001100000000010110101010110000111001100011111010111111011101011010101000111011000100000100110110000001001101000111111010011011100001101100110011101100101001000111011010101100010110001100110001011110100001011111111011010110001001011001000000000011000101010001101110010010010111011100010010111001101100001101111100110101101010101100010000110100100100101101010110000111101000000110001110110010011100011010001010010110101101001011010001110100110100001100100001111100111111000111011101010101110101111101011001110111011101001010111011100100011001100101111000010101100001010011000101001000001111011011101001011010010101111010101000101001000001000111110101110110011010011011000110000000011101011000001010011100001100010000010100111011000001100100011010110010100110101001110110001110110001000000100001111010101100010001011100001001001011111101110011001000000111101011101001000011001001000101100100100101000101001101101001000010100010010110100001111101100110100001000110011100001000101000000001100100000000010010000001101001110101001110000111110000001110010000010011110011110001101110000011011000110100010101111101101100001011011101100000001000110000010110100110010100100011001100011111000101000011100011010011111001111000111001100111000111010101111011110010010100000001000011101110010000010001110101111100010001110110001101000111100000110000000111110011001101010100111100011110111000010001010111010000111111111001001110101001010101000000010100011101010011001000011010011001011101011010011010010011100011001010010011111001001110011110111010000001100110001100101000111000011111110100001011111000100110010100111100010010001101010111011110000111000111011010011111111101010001010000110111111001111010001010001101101111000101100111010101100111100100111111100101111100010011011110100010100000001111000100011101101001010010111001010011110001011111101010001000100101110001011001000010100010010000111011100011010110010001000100110001100001101110000001011101111101010000011000101000000010011111001010101011101000001111011101111011011001101111111111101100011110101111100001001110001011101111001000101001001101110101101011110011111011110100010110000000101101101;
expected = 2759959;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);
#20;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd18;
noise_select = `BIG_N'b00100111001100010101010011111000010100001100110010100000111110011110100010001000100111000011010110001110100101111000110010100101010000111000111011111000010100110111001100110000000000110010010011000011110000110000010100001000110011011101010000000110101001110001101101001110111010000011011001101101110001011111011000111111011010011000110000111000111000110110101010000111101111011011101101011101011101110111010011100011100111001100001101010010110110111000100001101110110111111001011101000001000111110111001101100110100000101100000110101101111001100000000010000001001110011111011111001111010110110110000111011001010011100111001100000000011001101110010010010000000000111011101110110110111100001010011100100110011000100110101101010100001000101111111011101110110001011010010000001110100001101010011001101100011110010110000101111000010111110000111110011110001100000010000100101110111100010100010111100110010110001011001101101110101000001110011010000011101010110100111100110110000011011101001001111100100110000101000011111111001000110010000101110111101110000110111001000000000000100010010100011111010010011001111110000101001000011011100101100100100100010110010011111011010111110101110101001001001000101111010101111000100010010110101010101011100001011101111000111111101110011100110100001100100111111101000100100100111001011100100001010110011011010001001111010101111000011111111011111100101100111011000010110001111000010000001001110110100110101011110011101010111100011001010101100110001100100010110100101010011000100111101001001101010101001000000011101011001110111010111110110111110101101111010010011001000011110101011011000001100011000000111111001101001001101011100100111111010100100001111011000110001000001111001100110000111000110010100110000101000011111011010010101111001100110001001010000000011111001100010000011110111010000011110001010000010100010101001001001000000011101011110011011110000111000111010000100101000101111011001011001001001100101111111010111101111000101111001010010000011111100110000110011100110010010100010010111010010011000110000111100100010011100010100100000111000011111100010000001110010101111100011011111110110111101100100000101110111111011000000101111010100010000010111010010111101111010100001111100001011111001011001100000001101101000010000011000101101010001100010100110110001011100101010000000110011111110001000010110100100101010011001101110011110101110100000110100101111111001011000010000000001001001011000101100101110111011100001101101110101010111111110110111001001111000100110111110011101101000001010110011011100001000011111101011000111000110001111111111000111100000000101000101101001000110000111111110001111001001111010100001000010100010101000100100010110000110011011101110010111111000000011101001010011000000001010001101011011111001101011001011000010001011001101101100000101111110100111100000000011111011011100111110111011101010110100111011101110010000001110000110100011010011110001100011011010000011111010011010100011011100100111100011011111000001011111011010100111111000000000011111011100001001010100011100011111001111010111100001010101010101100001011110011100000111011010010001100010100000100001010111111101111101110100101110110001100010100011100001011000100111001101101100101000010010000010010101100001111101011100011000011101100001110001011100000110100101110100111111101001000101001101000100001111100011101101110001100011110100011110101001011111101010111101110111010111001010111100011100110011001100001110010000011111001111000111101100110110000010001010001010111010111100001111000011110000000101110011000101100100100100101101000111100010101010001010001010010100011111110100111101101000110110110000100101001001010010100011111001011000010000000010011110010001110111110100010101000101110101100110110111111110010111001100110110011011010001011010100001000000111111110111110010000101100010100100101001010011100110001110010000100110011001010101011001011111010100111101110101010111010010001101111010110110110110011111011111100010110100000111010011001110101110000011010101100001100011110111101001101111000101001000110110000101101110110100010001110110101001000111111100011011100101001101110000101110011110000100100010100001100101001001101000001011110010101011001000101100111100000111111000001101000010110000111100101111110100010000110110101011010100110111110001010111010100101011000010110100101011000011111101110100110000100110010011000010001010111100000101011110110110011001101000111001010100011110001100000100011001010000000000011110111001010000001011111001010100100000101000100010000100111010000110100010110001100011000110101000011110111100010010110000110100100001110110010111000111100001001001111001001001010011001011011011111101100110101001001100000011100010111110010111001000100010011100010001011111111011100110010101101101010000100100111001101101111110110101101110000101010000001110111011001000101110110101001110010110001010101011101100011101010011001010111111111111010011011111001100001010110001000001010010010101101001110001110001100000101011101100110011000110011101010001110111011100000010011100010110100110101000101100000101000001101111101101111010110000101010101001010101011111101111000001100111011001110010111111001011111001011111101111011010110010110110110100110010000010100100001000100000100101010001011000011101101001100100011001110101100001101001110110101000011111011111110010000010111000000100011110101111011111001011001001110110110111110110000011110000111100110101011001001111101011011000010001101110000000111001111001011101110000100010011110010000110110010001000101000001000010111010110011011011110000010110011100111010111111111001011110000100011001101001110111000101101111000101011101110011011100110101011010110100011110000101101101000100010111000000011101011111000011100010101011101100111000001111001101010101010100111111111100111110010001000100100111010010000111000111000000100011010100010110011111101100100001110110111010101000010100111100011101110000011011100111001010010010000101100001011110100001010100111011111100111001111001111110110001011111001011101011011001010110011100110000100111101100101001101100010111101000110001110001111111001000100111000011101010001011110100010110101100001000010100110010101001110010011010100110111101101101100010001011001110000011010100011111010010100101101010011000001010110100110010001000110001010010000000101111101110000110011110011111001010000010011001000111010000111111101101100101100000101110110010000101010010010111111110000000110010001100011100;
expected = 423326;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);
#20;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd19;
noise_select = `BIG_N'b00101111111000111110110000101001111011011111000000000110011110000001010101101001000111010011011111101111110110100100010010111101111100000111111011101101100001010101101111001000111101011000111011101101101011011101100000001000111110001010011000010111100111001111111110010100010100100000001011010000101001000110011000111011100100101011111011000101100000110011110101000111100111001011100100000010111100001100111000111100010110001011100011110111110011011001110110000011101011101010110011001101101101111001000110111011100000110000011110001111001011000011011011000101010001010111111000111100111110111001011110100101110100000110011111110110000100001010101010010101011100101011111111100111001110000110000101100110101001111100011001101011001100101010010111010011000101010011101000100010101110000100001010011100010001100011101101011011000111100101100001000100000101110001100000001110001100101011010110001000011011011010110011001010001011111001000110111010010101111100111100001110111010010100111111001011111001101001001001100010111011001100101111110101000111110011011100101101110001110110111011000100101101010100111111110111110010010100100101110010011111000100111100001011011000101101010111010100011100111110111011011111011010001010000111000111101011111011100100111000111011110010101110011010001001010011011010101101001110001100111100000000001011001110100001101111100100011100100101110010010001101000010110100011011000011110101100011011000101010101001111110000001011101001100110110101010001011011010101011001110001110101111100001010101100010111011101001010010100011100000110000111001101010011010100100000000011111111010101110101000001010110011101100010011101111000010010011111010101110111101001111001101011101110110010110101111110100110010000000110010101101001010000111011111011110100010011101101011111100100101010101111111010101011101001011011111001001001101100111101100110100111101010011011111001101100110001100001010000000010101011100011110101100100010111110010100101110000001000100110100011101110000001001110100101101111101001011011001000001110011111100010100110100011101011011101101101110001011001100111100111111000100101111000011000010100001111110001000100011010001100000001000111100001001000110000110001101011110101111010010011111100110010001111010000001100001111010100000000100010101010011011100011010001000000110001011110101100111001110110100001101100101111001110110000101111011000101001011100011011011111011001101011101000100111010110101010000101101100100101100101100010000011000100110001010001111100010101101111010101011100101000100010001110011100001111101000010011101011011001111001000101110101011110100000000000011101000000100101000010111001101110011100101100111000011101010001110100110101001001011111111000100101000110110010110001100000000000101011101100110111101111101001001000111100010001101011000101011111111010110001000100000110010110000100101111000110011010001110111010110011000100111010001001101111111111010101000110000001010001100010100101001001010001100100001000111101100010010100000111101111000111010000101101011011010110001111111100010000111010001111111001110111100001100001101000001000011011000100010110010100111011001100001011100110110110010111000100011110101101100001110001001000111000100101101001011111000111100101001111011000101010001101101000010100101101010011011101100111101001000001100001011101000011000111100000111111111100100001011010111011111110110000000111001000110101100010001100010011100101001011001011100000101011111000001000110100000110111110101010101000100101101100111001100111100110010010001110000000100010001100111100101101011111110111010111110111001000101110110110100000010000001001101001111111110001010111001010101100110010010010111100011101001111100000001111100001001110100011111010101011011010010001110110111111001101011111011110110110001110011010100101100101001111000011001101101000000110101111011101010001110101111100011101110100101010110111101110010110011000001100011000010101000110101001000111010010100011000100000000100101011101101110110010011010010100011011001011110110100100111010001000011010010011001111011000110001000001100110101110001000001000001110111011000000001010001011100001000111101111110000000011100101011101101010100110001100100001100011111101101111101001111001100011010011100011011110110111100101001100010001110101000101111010000010110111011000101110110001001000100011101001100001100000011000111110111100101001101110110101010010010000111001001100001100001010001100001000010100101101010101001001111111111010011000001011001011101100011000110001100001110011100010000010110000110100111010000100111110100010011010001100100011000111001100110001111110001110100110110000110111101001001110101101010110110001101111010110111110001100111100110101000110111101111111011001011011100010100100011010001110001010110111101010010111011100100111111011100111100100001100101010111010110000101101100011111000000000101000100000101001011001110011010010000011001100011011101010100010000110011011110011110001101010001111111111100101010010010010100000001111101011101110010111101010111110001110101100100001001111111101000100101100110110001101111100111100101101000011001110110110111010110110100010001101101110001100110011000101010111111011000001010001111000010011001011000010110100001110100011100100001011111110001101010110111100001100011100001001011111101000111011011010100000111100100100110111100001111001111010111110110000011011110111101000101001000000010010110001101001101000010101000011001101001010101111000111010001110000111001111010101110011001011011010011001010011111010100100010001010010011110001011011000110100011101111110000010101111101100011000111111101000000101011111011010100010100010000110011001101100000011010111110101000110101011000100001001011110111010100101011000001110101111001010101110100000111100100110111011010111110101000001111111101001110101100111110110011110111110100101110011101010001100010101001101001010110011000000101110101100011100000011011110101000111101010000011001111110110101001110000011100010000010011010110010010010100001100111001010000110101100001001110110110010101101001010110100101110100001111011110100011010000011100010000010000110011111000010001110001011000001111100100101010011100111010110011001011001011000001111101110000011110111001111010100101000100100101110011110010000101111000011101000011111010101010010111011111001001100001100101011011011111010001011011001001010010001100000001110101010000110100111000001001111110001110110110111001000001111000111001110;
expected = 10391768;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);
#20;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd20;
noise_select = `BIG_N'b11011010001111010111001101010101100111111100000011011100100010101101001111100010110111001100011100000101110101010110101010001111000011010111110011011000100001111101101110000111101100010010110010100101111000111010000111000000010101100100001110110101110010100010100010111111000001011011101100101101111010111110011101110110110100111101111100100001110100110111100100011000111001101010100010000001101100011011111101110110000100110101011000110111111010010001000101100000011110101000001100011100011110101001011110011011000100110110101000000000000111101010000011010000110001101110110000110110100010101110110010110101101000011100001001011000111100011011110011100110001111001100011001000011111001011110001101011000001111000111110110111100001010110110100101010101011101101000111010111111101000001101000010011110011011100110111101011011101101111011000000011100100010010101101000001110100101101111001101001111011111010110101100000000011100101111010001011000101000000101001101011001110100111101000111100010110100001101010011000110110001110000111101000011001111100101011100110001001001110110010111110100011101110101110100010001111001010110101101110100001100111010011111010011110010010000101100001001110010010100111001101101000111100011001101101110100011111100101000111111101011100001101011101111100110010000101011010100001111011110100110010001000110100110111010000000100110101010010001110110101110001001011010101101000011010110110101011011011110001101011011000101001010100101000011011101001101111001011011101111100100100110010111011110000110111101110100010000110000100001011000011011110111011010001101011100111101101111100101000111111000100100011010111000000110111010111010010010010011101110101000111101011101100001100111101101111111101101000011011011000011101000000110011001010010110110000011000001110100000011101001110110010010000111010000100000000000100110000110000011101001000010111001001111100010011001110111110110100010101010111000011110100001010000010011101011100010110000011110001001100011101111011010011011010111101111101011010011011000000000001111010010110011000111110011110000100101010100100110101010010000011110000010000100000011000110001110111100100100110010011111110110111111001100101000010000111100011001001111011100110011110010100011110100100000110010000110001100101010011001101111101000100101110001111100010000100010100000011011001000101100110110111010111010100001011010011110011100110101001101000110010111010011101000101010110111010101010100111101110000000011000011110000110001000011011010100111111001010100000110001000100101111110010010000111011100000110110110000101001011100000111111011100000001100111110110011001000100110011011100101001111110100000011011101001001011010010100100110111001001011010101001100100101101100100101001000100101100101111100101001011000100101010011101011111100101011110000100110101001000110110000010101001001000110001011101011000101100011100110001010111011010111011001110000011000000010000000111101000000110111100101001110111111010100000100001000111000111011101010001101010111010000110000101110010000011100110010011000011111001001000010000010001010110000010011101001100010101101011010011000100011110110001000001010110000100010010010001010011111101011001011111001010100010000011111010101110011111001100101010001011100110000010011000011101000000101011101011000001100010001110000101000111010111000111010000011010110011110001111000011011010110100000110000010111000010011000100001101010111001100000011110110100110111000111010011100011010000110110110000111100110100101011101010000100111100111010100010100111101100100011101110100100101110101111000101001110011110110101010011110011110101110001010100100101110100011011010001100011101011001110111011110011001100101000101110111001010101101101011000001001101101101001101100011101010101100011111100000110001101110100100011111101010110001001110100000110110110000000100011000101000111010000100101011111010010111000111000111111010001110101110001001111101100111100000001011000000001001110001101101000011101010001111010101000101111001011011101110000001101000101000101011110111010101110101100011001110001100000010111011101101001100100110110101101000111110011111010001110101100011000010100001100001111001001101000011111110001010000111000110101111001011111101010001111000111001101110000110100000110110100010000101001010010100110010100001001010110010101101010100101010101101110001101000101101010001101010000101011000011001001111001111101000110100100011011100000000111101011011011100110001101101001111100111110011111011011111110010001111110101001011101100000111111101011000010000001101011010001100110011100001111001011101100010101011010111101110100101011101011011001110111000111101110101011001010111111011001000110000011010000110000011111101111111111011010101110101110011000001100101010010001101010010101111111100011011100011010010010011001100111110001101100001101001111101111011111011101010100010100001011001110111100000011011101110010010011111111110011101101111000100000111000001111111011001100110100010111101101111111010101101000000100110100101110001011010010001000011111101100100001100110000011011000010110011110101000001111100101011011001100101100010111100100110011000010010011110100111111110100101001000000101111011010100110101110100001101100100011011011000001111100011100000111000110100100101011000111101110110111100010010100101110100000100011111100010011111111010011000100100100110101001110101001110010000111100010011010001000101001111001001111100111100111110011100010000010111001000010011110100010110010101001010001110010010011110110111010010110100010101000110011110110011011001101011111001010000010011010111101101011010010100110001001001101100010001001101101000101101011011001101111110101110011110101001000010010101000110011100111010101000011011000010011001011011000101110011011011001100111000110011001110110111000110111111011011001010011010010100000000110101001011111111101010101011010100110011000000000001101010000100011111001100101111001001110000010100101010100001010000000010001100011000100110000011001100111000011000001101111010000100111110110100010101110100010010011111100110000001011001101000000011001100000001111001111010111101011110000101101110011001000001011011111001000001111011100000110000110100100001011111010010010001110111001100110010000111001110100011101010011111010100101111110011110101001111111000111011000010111110001011010100100000101011101111100110111000001001101011100001010100100111101000010010010111001101111010010001101000011111111000;
expected = 9517808;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);
#20;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd21;
noise_select = `BIG_N'b00111000111100010110000000110101110000010010111111011001001110111010110110000111011001010110110100110100000010101000011110000100111001110011001111100100001100111111011101010010001010101110100010000001111111111011110100100001100000010011101111110110110001000011101101110011010100000011001000001011001000111010101110011000001101110001111111110110001010111101101100101011011011011111001010111010111110011111011110100010100000100010110001110101000111010001101100110011001000100000011010011000000111010010101110100011101010110010111000010111101010011000010101100011101111101110011110110100010011101101110100001011010000011111101001010000000111100010011111110000001111111100000001010001010000110111101110101100000100101110001111111011001011010010110110000111010011101010000010110101011110010001100101000011111001010110010011101010101011111000101001011001001100011011100001111101111111011111001101011101101110001110110010100100100010100011101101110111011010001000010111011110110001100011100000001000110100000101001110101101110000010111111111110011011111010101111000110101101100010001110011101101101111010001010010010110000110010111000111010010101001101111000001111010010010010100010111000011111001100101111100001010001100100111110111110111001110010000011000110110001110100100110000110011011011100101011000110000000010010011111000001010100010010011110100111110000011101011011000100011110011010111111001001101100111111000010101110111100111001000101100100000110010101100011111100010101001011110111111001101011111000001111111001101000101000011111101101101101010000011101001000111101101100000110110100110111101011110011000101110000100000001011101111111110100100111010001011000111100100011010101000010110010001000000010110100001110110100001101101100011011001110100100101000001111010110001111101110110101100111101000011111011101010001010101110011101001001100011001000100100011010001010000110011110110010000111111101100110001111101111100011001000011110010101010110101001111110111110101110100010111000111101101011011010111110110100100100100010011111001110011001000001010101100011100000111000010100101101110110011010011101111000101010001111010100001001101100101010111101101100011001111111010011110111010101000111100010100110101101011101011000110100001110111101010010101111100101111000010110010111111100111001110010111100000110001010010101011110100011111110101001100010111011111010100011110101000110100110011000110001101110110011001011011101011001110111001011000000101111110100000101001001010011001100100000011010111110100011101101111010010110100010110010001110010100111010000111101000001011101110000110001001000001001110111000100111000000010110011000101100111111010110010100001001110101111011001100101000110101100101101101011100100101111111111000000010111101101111101010111010100011011110011111001111000110111000000000100110101111010101010001111000000001010001000100011110001101110110110100101101111000010101100000101011100111000000010001111111111011010111010101100110010100000011011001001000011100100001010001001100000001101001000000011001001110000001000011110100100110110101110010001011001111101010101101111111110111100000001101011000101110001110000100001011000110011101001100011110110101010111001011001111011010001100000100111101101100101111100011110000111010001110000011001111010100110101111111000011100111100110100001010011101001001011010101011000100110011000101111111011011000011110110111010101111001001001100100100101010110001011101111011101011111111110100011011111000001000111110111011000101011011101011100011011001001101100011111101110000111010001000101000000111101111010011000010110110010110000101111101010010110011101010000011110101111000000100000111011001101111110111001111010110011010100010101010110011100111000101001110110010110010010111100011011101001111111011110110001110000010011100101110100100110001011000111001100110110010101001010101001000011100011110101011100000111011001100010011010101100101100010000110010001100001111001101100000101100000001010100010000101101100011011101010001110111011110111001000101001010010000011111001111010011001101011101001100010110011000000111110100010011111110100001111000010011101101011000110010010100001001111000101011000010100010000101011110010111001110110011001000001011010111101100001011110010010101000100100001101001101100111001110010101000101000111001110100000101100001101100001001110010010001011000110010000001000110010100011111010110101100001101110011111001001110100110000010010111100001000101101000001111100011000110100110001001100101111100100101101011011100010100100110010011010111100011110000100100101000110000010001001011011000101110010100011100010010010111001110110101011100110111000100001110110001010010011101101010101111111001001000011111010001111010111111110011111010000100110111001100101010011101011000011001000110100000010000100001001000001001011011000011011011100110101011110001111010010010100000111111011010101011001010000101111010011011100010111111111100111000011000100001100011010000110001110000101100011101111110010100000100110000100110100010011001011001101011101110001111100101001001111010010001010100101000000010101000101011010010011111010011011000011011000100101001000101011100101000000001101110010011010111100000010100010101110111001110011001100010011011010001100101000001101111110111101010010000010010010010101100001110100111110111100100100101010111001010010100000011000010001101000011111001010111110100101010010000010001101011100000101100011111010101100010000011101000100010110111100101011011011100101110000101010011000100110100000010111111011001011101111101110101010100011010101010111001111001101001101011011110111101110011110010110010010001100101100110101110111000011000111010110100010110010100001100010101100000110100110110111110101011001100011000011110110111011100100001101011000010110110100101000111001001101101101100010010011011101001011110101011111110001110100000001001010011001001011000110000011101010100100001001110010101100100000000010001001011010010110001111010011011100010111101010110000010000110000010000001001000101001011010000110110100000011011001111011100010001100100000111001111010001111101110011111001000101000000001111101101001110111001010110101011001101011111001111000111010110111100011011101010011001001011100100100011100101100001011111100100110110001011100010110001111110001110110100000110001000111010100011101111000111011111111100011001011000100100011010101101101100001100111001011100101101001111111101111011011010011011011100011101110110100;
expected = 9315338;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);
#20;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd22;
noise_select = `BIG_N'b11100001010011011100101101000010101101110000100011000100111111001111111000000101011011110101100111001111001000110110011000111110001111100110011111011000100001010110011111100011100000101001000000111101100111001011101001110011010110010111001001011001011010011010001010010010010011001000110011001110000001011111000011000001111001101110011101001110001111110000011000001101100010111000000001110001100110001010001011100011011111111010000000100101000001101001100111111000000111100101011001000010100011011011001001010100110101110011010111101011110101100001101101100110011000110111001110111011001100000110111100111011000100101011110101010010001001100100100010100010000100110000110110110001000111010110110010101100011001111111000001000110001110100001011101101001000111010000100100100110011011111000010110010100100010011011100010001110000011111101010111111111111101010001001111001011011110011001110010100010110101111011000011001101000101001110110000100101100111111001111000000100101011001111011000110011000000010100100010110011100011010011000111110011110011101101110111000000111000111101000111000011100000100010101101110100000100101011101110100000101111100111000000010001010000010010010011010110010010100001000000110011111000111100011010111111101101100011101011001110100001111001111110010001100100100110101100110101011011000101100111110001011010110101101110101000001110111101111111111100111011110111000100000001110001001111111001000010101110100101111001100010000111010001000110100100110010100111011111011111010110000110010010011111111101100111100001001101000100110100111101100101010011101100101111001100000101000100001110001100110111011101010110000110000000110100011100100111100101011110011011111000001010011110110001010110001100001111111010000110011011101011000011000000011110011111011110010111101110001110000100111001100011110100111010000111101111101100010010110111000101000000010110111001101011100010101010111110010100010010100111111000111110100001101111010011010111000000001100000101111000101100011001110100101000010100110000001111101111011010010000111110110100001011000010101111111111100011100011011001010011110010000011010000110111001001101101111001001111010101011000001100110000111001100100010110110001000111101110101001110011011000110000100011001110101100111001001001001111011100011111010001110011111100100000101100001010101111000000011101010001100101110001000111110100111100101100111011100100000111011110100100010100000101111000011100001001101010011111011110000110110010101001110001001010010010110011011001000100011000110100100010100010101000101101010111001001110011101100011100101110101010010100111000001010000000000001000111000100101100100111111010111001100011100100001010011010101001001000100101011100001101011110110111101011110111101100000000010000110001011110110001010110100111110101100111101100010100001010000011010100001100000001101001010001111010110010001101100011010001110000111111010111110001100110100000100110101001001110001111011111000100100110100101110000100011100010110110110100010010100011110100011110000101111110001111101111011010011011100011010111110111111100101010000001000100000101100111111110100100110110100010011101010010001010110101011100011010100110100000011000100011011110001011000001101101100110111111100100011010011110000101101001100110111011111000011111111001100010010111110010101101101011100100000001110101000101110111111001101010100101000011010011010100001010011000110100001011110101001011100110010111010010100100100011110010011001110110110001100000001010100011011110011110101011101010110010111101011101100011001101001110100000010111100101111001010001111110110110111010010011101011000001000000011010000100110111100011100010110111110001110000110001111001111010111111101101100110100011110011000011000010100101001100111011101101011100110100011000001111010000000101001011101011100000001110001010101010010110001000000101111010110101100110000011110100000011100110001110000001001010100101000110100111111001001001000001000000000111101100111101100111000101000010001010110000001011001101111001100010100110111100010100110100000111000000011100011010010011001100011101101101000001001010111110100010010101110001101011111110101011010110100001101011000101100110010111000000111110000110110100010101011110110011100010010001101000101000011110101110100111001111011100111001001011100111001111101111100110010100001111111110000001110000110001100011110101001000001010010010100100110010100111101011011110111101011110101010100001001000000111011010010010100110000000111000000110010111000001111001100000110101001000001011001000111101011111111001010001001010110101110011001101110000011001010110001101100110110000001111111111100011000110010110010110000011111100110000100011111100100110001110010111100111100100101100100010111001111111011011010010001100110100100110001000011100110111010011100111110101001100101110101000110010001111111110100101100011011011011100010111110111101000001010111001110101111001010011000000110111001001001100001101110110100111001101010100010011111010011010101110101010111111110010000111111001110101001000011000010010110001110111110001110000111001011111111000000100110111111111111110010111001100111110001010011000011010110100001111111100001110100110100111011100110000110111101001010010101001010101010011010010100111101101100100101001101111111101111001111110111100011010101001100000111101010011010101111000001011110001010001001001011101110110100101110101010000110010111110011001111011001001011010100010101111110001010010100000010011000000111010110111101101100110010011101011001011001100010111100100100110100100010101010111000101011000000010011111110110010010111010110100001100011111001001010010010010111110111001000010000111110010101110010011010001011111011001111111100011100011100000100111100000000010010010000000101010110101001110000101011101110100011000010110110010011100110101001000000111101100101110100111010000000111000010011001101010000111001110111011000000010011100001010110001111011011110110010111111101010010101101110100001110110111100100101001011000100000010101100111100111101010110101110110110111110011010110111101101010000010110000001010100110011000010101110111000010101010010111101000001111000001110001110100100110101110000101101010010111100010011101000111110011011100101111011000011011111010111111111010011110011011111001111110100101111111000011101011100011000000001101010110010101000010111011111111110101011001000111100001001101000001011110010100010001000111000110010001001101101001011001111;
expected = 102016;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);
#20;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd23;
noise_select = `BIG_N'b11100100010011000100010010011001011101010100111111110001110111001100101001011110111010001001001101110000001000000110110110100111000101010111101111110001110000100010000000011000101000010110100101001010000001001001000010100111001011010111100001101110111011111101100110110010100101000001110011100111111000111011000111001101100001011100111000100001001001001111011000111110010010100011110011111011001011100011000100010000110011001111111000000000011001111111000110110010100110001011100010110110011101000100101101011010110111011000100000001100100100011001101110111011001101000100010000001110001101111011000011110000001000010100100011101101101111100100101001101011111010010001000000111110001111001010011011100000001100101101101101001100100100101000010100100110110000101100000100000000111111011000100100000011110000001001111001101101110011100000011000000110011111011001110011111100000110011011001110000111101111010010101100011011011110011110100000000010101110100001011101100011111111010001111101000111001110011110010000001010110001010110110001110001101111101011001010111011000100111110110010101101100101110010001101111101000010010100110110000001010110111110011001110000110110011001101110101001111010000001111110101101010111001101101010101010100101000111010000000001111101100100010101100010000011100001011110111100010111100110011001010111111011001100100001100000101111001111010101010100101110011101110101111000110000001101000001110011101101010000110000110100110111000011000101011100110100110110010110101111000001100001110011111001111111001000000111100010111100110000101011111110111111000001100010010110100110010001010111010101001000001010100001101011111001010011101010101110100101000011111000100010001100000111010111001010110010011110011001000011001110011101000110100000101101111100100101000010111100110101100010010101001111110101111100011010100100001001100000001100001000010011000011011110100101000101011111101011101100001101101100111010100000001011011110010101111010101101101001011110011100101101000111110111110111010000010010000000100011011011000111010110101110011010101001010001101110110111000110110111011101010101100000000110000100110010110101100111101110011111101111011101011000011101001011010011001101101100011011101001000010101011111101101000110001010000011100011011101111001101000010101000010111101000101100000100011010001011111001101111011011001010000111111101000101111001110101101000100110100001001100011111011110111010110000111000100000001001000000101110001100110101101110001000110110100111011100011110101111101000101110101111010111001010101000101000001111100110000111101010111101101010011110010011001011000110101100011010010010111001111110100000110100110100011110111000111001100110011001001010001011110100010001111101110001001110110010110011001111101110010111000100000011001010110000010101100110001100000001101000100110001101100101001000011001000000000010101101001011001000110001110001101011110010111000110010111001101001111111101000001100001110101100011100110000100100111001000111111010011001001010101010100010111010000011011110101111100001100101000011001011010101010110010010110000001101010000000011110110011000000010011011111011001110010011101000000110011001100000000100110100101001111000001010110110011101101001111000101100001001100100000111110000111010011111101100011001011101010001110101011100011011011000110010000101001100001010101000100111011100111011100111101100101101010101001011101011100100110000100110001010011110110110101001001001010001100000101001010001111101011100001111001000011101010001100110000110111000001000100110001010100001000110001101110101001011100111010111101101010010101000001101111100010110010001010100011000110011110111001000010000100110101111001000111111001110010110011110010111000000101001011101011100010011100001110011101111001010001110011010000110111001101000110011101011100110100010110010100110110000001101101100111001111110011100000001101001001101111010110011110001010011111101100000010111011000010000100001101110011111010010100100010100010111110001001000110110110101010001011001000001011001000110011000011000010111000110110101010010001001011100100110110000100110000011010111011111111010101100010011011110010101100111000101111100110010111001000111101111000100111100100011101110010001111010000111010100011001001000110110111110100000010100000111000101111010101100000000111110100101000111110100100111011101011011010000001011011011010111110110001011111011100110010001000001101001111100111110010110111010000000110100001011000101100001101101011010001111001000001101001001010110010101100010110010110110110110101011000001010101010100001000100001010010111001110001111110101110110101100110001001100010010111001010100010000110100001010110011110101110001001000101110101110010000110010100001101111000111010110001100001100010000010100110110111101100010001000000011000001101000110010001110100011111111011010000010000000001010010100111001010111011010101111001100011110000100110111110010111011101000110001100000111001111010010000001000100010011010111000010110111011001110001000100101000000001111100111001101110000101110010011111101101001000111111100101011100100111011001000011001111101100101001101110100110101001001111100110010010010100000100010001111001100101101110010100001111100110111000011110001101111101010010111111100110101100010101111001000100011011101000111011001101011001000001000001000111001100001111110100000001100111001101101000000001001000101111000010101111000000110101101001001100001101111100111001000111110110011100100101101100001110000011010000101101111100110101110001001000001011001010000101100011101011011001011100100000010111110111100010001010111000101001101101011000011011011101110010010100101100001000000001010111011100010100101011010010000110011000001001110101111000000001111000110101111111011010000000111010010001100111010110101110001000010001001101111010100110011110011101100011001110000111110111100010111111100110011111101101010111010011011110000111110000000010111110101010001000110111111001010001011110111010001001100100001010011101111100100111100111001001010001111111010101001010001001010001101010101001000100101000100001111010001101110001011001010110011111000100100110010001001111000111110010111110001001001100111111111111010100110100110100011100110100000010100100110010000000100100100011110001101010101111111000110101001010110010111110000110110010111001110101101001000110010010010110101000011001000000010010011010011001000101001010001111000010100000000001001010010110110100001;
expected = 6407664;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);
#20;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd24;
noise_select = `BIG_N'b11010111100101001101111001101000011001110110111101111010101100010000100100000101100010010101100110111010011111110110010111111100100011111111000000001110010000011100011010101110111010000110111100011101101111000001010101110001100101101110110011001111011111100010011111001111000100100100001110101001001111110011111011101000000100101101100110000101100101111010000111111010001001011111111111101000101000001010000110010001000000001011000111101000110110111111110010110100111110011000100001011010111001101010010110000011000100000000000100101000100101110101111010000001000011000000001001111011100110010010001101000011110000100000101111110001110000111001101000111011011000000000101000000011000010110000001110110100001100111111011100001011110101100110011101000000110010001011101011100001111101110100011101011000101010011100111100010000101010011100011000101110011111011011000110001011111001110001110010100010010011000011011100111100000111001001010001011111101010100000111011111100100100010111110110011101010010011111001101011011001110100000110101001100001101000100000010110001111100111101100010000000010100101111000010110101000100101011100010100001100011011110010011000010010111011110100011010100011000111111001000100101001110011101001010110100000011000001011001000100110110111001101000110010000110010010000010001110000001101100100011100110011101011000111101011101001010101101100001111111101001000111000100010001101110111000000011101000010111001111000101111000011111000001100001000000110110010110111010010001001110101010110011101100101101000010001110100111111100100011011000101010010110111001011011010000011100001000110010000101101110000001111100001110010011010101010101100000111110111011011100110101000001000011011101001100111011001011001101100110100110110011111110110100101111100001000000001001111000101111100001011101001111110111101101101000101001110101011011110001000110010001110111101100110010000011000110110001001001001101000001111111011011101010101000110111100111000001110011101110000010100001110111000101001010110001101111000111001111100101100001100111111010000100110010101010010011110000111100111011110011110010011000100010000010100001100100011110100001011000011011010011100011000110000111001000101101011010101011110001011000001010101111001010100101010010011001000010011000001100010001100110101001100101111010001111000011101000110100001100101001110010111000000110100101100111011100000011100001110000110000101000001000001011001110000111001011100010000110111011000011011011011001100000101100110101000011010000111111000100111100101000000101001000011101001110100110100101010010010010111110100001111110010010100110010100100010001110101001111100011011101111010001010111110000011010011000111110110011110100101001001101001100000000100010010000001010000101101000101001110011010110101010000000001010000101011100100001001011001101101100110001011101110111100000111110000101100100101011100111001110001100101001000100101100001000101001110111011010001011001011011010111110000101100111000101001110011001100001111100000101100000001100000000111101111111011110011010101100000100110010110101001001101110111001110100000010111001010111111101100101000111110011100110001110001010001010001101000111010110001010001011010111101110001011111011000001101111001001010110000011110010011001111001011111111111111101100001111011111011101111001101001110001011100001110010000111011100010101110101101001111000001110111100101100010101111000110010110110010100111110010111011001111101100010000011101100111101010100110110011001011110100101111001111100110001001010101100100011001100000101111111001101000111101001111110100110111010110101001100010000111100100100101001001101000001000110011011110100011100100100010101110010000001100111101101111001101011000110010111101100011100100101111000010011111101100001010000110011010000101101110100100101101001100011010001101100001011010011010010111110111110010011000101100100100110010110101100110111001111001101101111011011001010100000101111100110111100000010110001111101100000111110100001000010111001111000010010001010110101011100100001001011010100110100001001011011000110100101110100100001001110001011010110100101000010011110100001110110111000111111000100000001101110001100001001101101001001011100100010000110100001011101000001110011100110110000000111011001111111001111110000101011010000011100111001101101000111100000100101010011110010101101011101001001110001011101000001011011001001111100111110001110111010011100001111101110010000000100101010100100001111011000100000101101010110000110100001011001101110001001000110111000000001101100100110101001100101101011000100001100100001010001000110101111000111100100001010111111010000010111101000001111110000110001111101100111010110111010000001101011101100001001010011011000110001110101011001001110110001010101111100011111111111111101001111100011110010000000001101101101110111001110111010001111001010100011101011011100010011000101001100111101110100110110100011101101110110101100000000111111001101000011010001001100001100001010111100100110000001011101110001100010100000100000100011111001111110001110010011010000000111011011110001110011010100110110000101001100001010100010100001011110110100100110000100000010110101000101011001101000000111111011011100110000101100110110111110010011011001110011010001110110101000010101110101100100011001011011110100010111000100000100010100000111000011110101001000110111011001101101100110111100111001110000011001111000001100100001110111011010101010110110110100101111011110010101011110111110011101111000001110110101010101001101111011110010010001000110111001110110001100101011010100001101001011100011100010010100111101100010010100110010110101111110011110011011000100011000011001000111110001110001010000110011101011110101111111011110010111010100000010101001011010100111100010010000100110000011000011101000100110000110011111010001000101010111110010001100010111100001100101000011000111011100010110001000010110110000010110010001111101110110001010110010000000011011001110101100011101111000111100100110010101101001111111100001010110101011001110100100011011100101000001100111101000001110111011001010110101111110111101101101101000011010111101001111000100001111101011001010001101100011000101100100101001100100100010001111110001010111011011110101010100001111010000010010011011001000001111011101110111000101011111111000001101101011100011001010010001000010011100010101001101001110101101011100000000011111101100100001001111000000100010110110001000010111101011111101101110010100100;
expected = 9729564;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);
#20;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd25;
noise_select = `BIG_N'b10111101000111011111100010100110100110010100110011101100001101101000011010100111000011010101011110110100010101101001010011100001011100000100011100111001011001100101110101001011100111100000011000001000001011000001001010011110000001010010110100000101011000110010111101010111101111111000100110010100100111011111000011000100110100001001011011100010111001110110100101101000101000001100000110001000110111101011101110101010010110111110011000010100000011101010100101001011011011010011011101100000011110000001111111010111001000000101010101000101011001101000001011100001010001001000011011101011101111000100010101111010101101001001011111101000000010011101100011010111111000111101110011110000101010111010011000110101110110000010111000100101001000100101001101010011111110111111000011001101011010110101110010100100011101111101010110110011001111100111010101010010010011101101010111110010101100110110011000111000000111100100011110011100110001110111100000110110111000100110110100111000101011100001010110011101111011010011000110101111011110110010001110101001001101101110011001101100001010111001010001100100101001100000100011000010000111100011001010110100011111000000001100010010100111110001101110000110001011111000001101100110000111010111100100111101010001111111001100101001010110101000000110010011011101111001101011000110010100110100011100101100101101000010111001110110011100011001000000011010100010011110011101100000110111001011001110111111101111011001100110000001010001000110101011011100011010101001001110101101101011000101110001011110010111010011000111110101000000001011001110010001100100111001000011110101000111100110000110010010010000100001010000001100110101110001000100010001010011100011010011111100100001111100101001010101101011000010110011111010110101101001101100010001111101101110011001100110011010101011110100111011100011010011000010110111000001010100010001001111100011100100011011101101111100100010010110000110101001000111010000011110110001000111010010010100110010010000000100010101011000001000000000001001110111110001011001001110011111101100100100000001110101110100011100101100001000010100111100010111001110011111011001100001101001111001110001110010111010011001011011011110101011000000110111001010101110011000100100001101101111100100101001100100011111010101101110110001000111011110011101110101110001010011010000010001011000011111011010000110101101011010001110110010101100100100100101100110111100110011100011010110010000011010000011101110000100001111010100101001001000110110000010000011000000010101001001111000101000110101110001110000001001001011101101000100011101110111100010011101001100100101011000110111110001011000001100111110111110111110110100111100000111000001010000110001101011010001010011001111100110011111011110111011111111000110110101010111011100000100100001011110010111101110101110111111000100000010000010000001101101011001111011101011111100100001010110101110010011000011101100111110100101101100000100101111111011011001001100001011001100011110011000011001010011011100010100010010100010010000110110011010011010101100011100100000111011010100010000010000001010011101011010001011011110011100001100100111101101011100100101111101110010011001000010010100110000111011110100111010011000111011111101000001110101001000100000000010000001010001100110001100110001010011010010000101001000110010010000111010111101100010010100111000001110011001101101001110010001100111010000010011100110110100111000110000110011111101010111100100000011100110100011001110011111010111001001000011100110101110101010001111111001100100101100110000010011111010010111011011001001001000001011100001101100100111111110001100100101001111010101101010101110011100001111101001101011111001011111111010110110011001110011110101101101111111101000111001101100110011001110010100001111000110110010010110010111000100001101010001000101011100110100011000101001101101001100100111100100101000111101100101100001010100100110010101110110101100100010000001010001001000011111010111110111011010001111001000001000010001000011110010010110001001010101010110010110111001110100000001000001100011010100110011101100101011001001111101100110101011110111010100100100111101110111111111100000011011010110110101100101001100110111010000001000001101011001010000110001010001000001001011000111011101110010110001110011101111100111110110111100110100000011110011000110010111100110110011101001010000010011101111111001110010111010101110011001110111100110101101101100010000010000011010000110101110001000110001110000100100010000001000101000001100111001110001101101010110001110000100010111100011111100010011111100110000100000111101111100001101000100100001110001111100100010000000000111001011101100111000011111001011110001110010100010101000101101000111011101000100101001100011010010111101011010111010100100010101111100110011011000100010111000110010001111010000011010011011000001101110110110110101110000011110101001101101110101101011111110000101101110100001000111101110010001011101111110100001010001001011010011001001010001100101001110111000001101101011011110000011111010110000011101011011010100100001000100010100000100010111011100001111010111111000011011000010011010010001000001000111110000110000100001010011101001101011000011010011010101110110111010000101100011110000010101111101111011111110100010011001000110100001011010101000100001000000110110100110000000010111101101011010000001001110011000111011000111111101110001010100111010100001000000000110110010100101001010001010100101100110101011010010000111110010010010011001001100011000111000010010110101010101000111101110011000100010101000001111100110111000110011101111101110111001101000011010110011001000111110101001011000111100110101010001010000101110111110001000111111001010000100110000110110100110101101101111111001110101111010101011001100010110101111000011111110011101000100000101111001110101001100010001100101001101110001001000011010001000100010001000011000010100111101001111110011111111111110101000000100010100000010010100101100111111000111100100000101100111111101100101110000000110101011101101110101111100010001001100101000110111000110000010010100101010100000001000010001010001001001110001101111000111100000000001000110101111101001101001001111001011110001011001101011010000010101111101000000010110110011000000001000000101001110110100001110111000000100010010101001011101110001100101001111001000111101000011000101100001011000001101111011111000111011111101111010011111000010111011000000110001011111011001111010001011010011110000001100110110110000110000100001110;
expected = 2066905;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);
#20;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd26;
noise_select = `BIG_N'b11101111000111010010100010010111101001111100111100000100000100111010100000101010001000001100100001001111110010001010111111111011010101011101101011001101100011000100011010101001011110000101101100110110011110101100101101000000111101100110000000100100000010001100110010110111100110101110001011001111010110101100010110011001010011010101010101000010010001010100000011110110100010001110111110011010000010011010111000110010100010100110010111000001101111011011000000010100001110100011011111111101001111011011000100100011110001101110011000011100100000110110010001001111110100101001011011001011011101101111111011100000000001111010100001101000110010001110010110000011011000000111011111011111000101000111001011111100000011000011101111001010100011001100111010110010111010111011011001010011101000000011110110111001110001011111001010111101101010010010111110100101100100111111000001010110010001110011000110011000011101110110101010000001001110000111001101010010111101100011101100100101010101100111000000110100010100010111011111110011111010011111001010010110001011000101010000100111010001000011111111101000011111100101011010000110100111100011111010110000001111000011100111101001100000111100011000100000100000100111011110110011111110100111010001010000011011001101100110101101101001010000001001000110101100010000101001001010001101110101111100111111010010000010011011100101001111011000100101010101101011000111101100110000001101001011111000110111001011011010111011110111011101111001001000101101110110000000101000100001111001010000010011000011011100001010010110101000001101001010101011100101100000100000111111100101011111011101000111001110010100110100001000001110010011001010101100111010000000111000100010000001100110010110111011000010001011000001011011100000001100000111110111100110101111100011100010001010010010101101000001111000111001100000001010100101101100001111000000110001000111100101111111011011110111011000110010000000000010100110110100011100101101010000111111011000011110110000011011110100011011101000011010011110001001100010111101101010011101001100111101100011101001001001110111100010001111111110110010110010000111100111000101101101001100010101111111001111111011000100010010101001111011000110110101011111110010011111110010111111010000111101110111100110011011000001111111010010100100100101010001100000011011101101001001101100101011100100001111011101110110001111100101010010001100011111001110110110011110010010101110011001011000111111101001111001111011111100100111100001010000111100110101110000110011011101111111010000111001001110011000100111001010100101000001111101010101101110001000010001010001010011011111110001111001000001100111011001001101001110010000101001000001100010011110000110001110101101010100010011000100110100001011010111010100111010100100010110100111111011001110001000010010010111010000000110001010111100100010000100001100100110011101001110010001110001110001001100001100110010001101100110010000001110101110010001010010011101111100110001010001110111011010111101111111100010110011000111111110000110111100111111111010100101000010011001111110010101111010100101011100110011010011000111011100010001000110001111100011110000100101001101111010101001101010111001010000100101101110110101000110011010110100110100000010001010010001001001001111100101010100110110111110111010010110011110001010111111000111000101010110011001101111011101000101010010010101101000001011111110100010011000101001100100111111011010111001111110010000011011101001000000111000110111001100000001110100111101111101100010010111010001011101011000000001101110000110100110011110001000101110111101000100010110101111111011101000010011001100011111100110100110010000001110100101011010100111011010010011010100001101001000110010101010100000110001010110110010000011001010101100110110110010110100001011100011100100111000001111000011101010010011100001101111010000001000001100011000101101101101010000000010100100110101000000001110010011110101000101010101010000100011110001101111001010110011001111111010001000010110111011111010101011011111001000101001011000011110100000011000011110010001010000000011110010011000001011110000000110011011100010000010100101111101010110101001110010101111011100101111001011000000100001011010011101101000001011101010100100111001010100110010011100100000010110000011010111001101001111110101101101111000001011001101010011111010100010100010010011011100110001101100110001001100001111011011000000010110001100110110010001001111001011010010111110001010100111000001100110100001101100001111000111111001111000101110011001111010101010101100111111100110101001101001000110110011011001110001111101011011110000011101110000011010011000010011010111110010111111000111101010010110000111100010000110011000100000110000111111010011011100000000101111100010011110011010101101011101010011100010111011100001001001000001100110000110001100100101010100111011011000110100000000011111100000101101011000110101100101000111011000000100010110010100010011011101100100011010001010000101100001110110011101100010100001100111110010010111001100110011011101100010011100011001001101001111010001000011010011010110011001110100010100111111010101001110010111101000110100001011011100100001000110001011001010000111100110111001101010100011100110100110111101101101000111100000010000000100001010000011110010001101110110011111000110100100011101001000110011111010100000100100111110111111111010000110011110010101001000101111000000111011001010000010000110011100010010111101000110100000011111111100000011001110110010110101000011101110100110101110100100000111101000100101011110001010101010011011101000111000001011111011110101011100100000111101000111100100001111100111001101001011001001110011010001000100011111100100000010010010010011001111100010110000110101011000111111011101010100100110001110110111010101110000100001000101011000100001000111101001101000001011001001111000001001101011101100011010011010110011001010100011110000101010111001010111000001110001101011000110111001101000000101001011110100110100110100010111100010011001111011000000100011101110011011101001001101111100101100110111010110000001110101011100001111000100100001111000010101010011101111101011110010011010100101101011011110110001110010101001001101000111100110101111110101011100100011101000000100010001100101101111011100011100110110011001111000111111001101111100001000010111000010000001100010100011011111000001110100100001001110100111010001110100101110111001111100001100111111011100111010101111110011111110111000001001001110010111001110001001101100010;
expected = 4524496;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);
#20;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd27;
noise_select = `BIG_N'b00000100111101110001001001010010110010101001001111011101111111101000010001101001111010100000000111111101011111111101110101010010100101001000001011101110001110111110101111111101001100101010111101010101101101100101101000101000010011111110101110101000011111001011101001001000100001000110101111011101011100101100101101010011011010010110101010100111101111101101101011001100100000010011111000001111111101001000110000111110000101100101101000111001101100100110010000011011100001000110010101111000011100110000001000000011000011011011010100000010100100011011101010000111000011010100100100010010100101000111100001000011000101001111111101011101110010011001101011100101010011101010000010100001000010000101100010111011101000000101001101011111011100101001100101111100110011011000111001001100101111011010000101001011111010100110110111010110010111101010100110100011011111101110101000111001010111010010110100111101110010001110010101010110111111111010000000000010101010010000110110000111110111101100000001011111001001010110101111000101111010010011110111000011011110010001101111000001100001101101011011011001111011101100100000000111000000111100001110110001100011011110001100001100000100110110111010100110011011100010010101111010011111111001110101001110001011010100101010101111000010010100111110100110010111011100010101101001101100011111000011101110101010001110010001101110111011101001110010110111011010111111011011111110111001011110110111010010001001100010011101010100110001011110100000100101001100110101011101101000100100101110111101111111111101111011111110011100110000101101101100100110110110100111100111001011001001101011111110101010111011010110011101100101111011101011001010010101011101000010100101000010100011000000111101100010110101110001000011100100011011100001010011100111100110101011100100111011110111010001100100111100100011101111100110001010110101110101110111111100101011101101001111111001001101110001001110001101100100100110110011100111111001010000000011011010011010001000010110011110001110011000010011010111111111110111100100111011100000110010101110010110100100111010110110000010111001001010110001001111010100101000101011101001011100001111011011101000101000111000001101000010100100011011000001011100101010101010011010110111010001110101011001010010111110010010001011000010111001010011000000000011011001001010110100010111101000010000110110111000110111100011011111001111011110011000110010111101011010001100011011111101111001000011101011111111101101001011111101011000111110000101001000100111001010010011011000010011100111000001100101101000100111010100111111101111000111110011101101100110000011101000101110111101000000001110100111111100001000111110011111010000011111000001010111011000010101001100100010110110010111101010011101101010000100101010000000010111100111000110010011110011100010001111000110000011111001100010001101101001111001111000010000111011110000100101010111010011010000001110101100000100011110111000010010110010101010110010101011001111011011001110010000110100101001000000010011111001010001000011011011001111010101010001100000101000111000110110011011100110000111101010110110111001100100000001111011001101001110110111000000101000001110100011001010101110011100110010111010000011010001010011111100101011101001011100101101000000110001001010000111000111000010011110001111000111111011000101101100110110011000101001010111000000011001000101111010111101101001000011001001000100111111100100000000011010110111100001111111011001010001110010100000000111111100110110010011111110010100011000000001011000010010101011100011101101101011010001011100110000111000111011011101110111101000111111001110110010100010001001111001111101100111101111100001010100011110100110001110010011010101000000001010010111100011001000010000011010011011101001000100101010100010011001001111111100001110011101111101110101000001001110010100011011110110011011111010001011011010111100110100001010101100011010000011111110100011110010010111001111101010111011010000001001110100011000101101010000010001011110101101110010110111101101001011101100011001010001101000100111011001011110001110110011001010100100001101110101111010101110111101011010011111000100000000001010111001010101111010011110110100000011111010001111010001001101010001011101111010010101011110000010010110001111111101000001011111111001010001001101101101001111101001011110000010111111111110001000100001010111010100111001110111010101001111000111111011111001011000000100001111010100110011111011000001011001010010111000000011110001111101010001111111110001011100000000000010000111000101111001011010110101000101101110110011111000000100011011011111001100101111111001110011110110100000111001010100100111111110011100010101100011001011111000111111000000100011100011000101010101111101001110001001101100101000110101111001010001101011101111001011001000111111001001000011001110000000111110011110101101000001001100100100111100100111101100100011011000101011001111100110001100001000011011001000101010111001000111000001000111111101100000101011000001111101101111010100000010111011001100011010100101000010011101000110000001110010000000011100011001000011000101010001101010111100011110110110000011010110100100000110010000101101011110100010101000000111001011011001000101101010100111000000101010110000010100000011000001110110010000111101111100101010001110011001111001110011100000011000001011100111100111101110001110111101100000010010001010000100111101101001100001100100011001011011000001101101000010100101011100110001110100100011011110111100000010110101111000110100011000010000010100000011000110011100001111011000100011010101011111100001010011100110010011010110010000110000110000100011010110111100110110010110001101110011010111000110001000001101000110001110010000100100101000111101100000000111100001000101011100111010010011000011000100111111100101100000000011111001010010110000011100011000111110010100100101010000100111010110111000001100000100011011110000000010000001110111010101010110000101011100011100010100101001010111111110110111011101011110010100010101011110010111001001000001111011011011001101001001111011011110111101111010001111011000100000110010010110000110110110011100010100010111011011001010011001001110010101010000100001100100100100010110011100110001100001101111101010111111001001101011011101110000101001011011000100010000000100000011111011011111010110101001111011111001011011001101101001011100000101011101110001101010100011010001111010110010010001011110011000101000100111100110110111001101000100111110000111101000011111110110010;
expected = 10913504;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);
#20;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd28;
noise_select = `BIG_N'b11101101110110001010011100001100111111110111010100011101111111011010010101011100101111110100010001101100101110100010101100101000001000111101111000110011110010110011000111101100010110101111100010000001011100010010100010001110110110101010101000010110000010001111001110010001001100010001000100001001111110010111011110111100110011100111000111101010010000101000101000111011110100110010111111100111010110100010001001001110110000010101101100100110010000110000011011111000001001111001111010010011011100100011110111101111101100010010110111010011011100010110010011111101100110010100010001101111110100100011010100101001001110000010110000011111110000100101011001111110010101111100011101011011011111111111101110101101001001000011100000100110100010001100010010110100110110110110000110100001100010011100111110101110001000101001011000011110110010001010110111011010011110111101100111011000000001101101001101111111111010110010011010111011000100001000110000001100111011011011100000111110010110111001101001010111111001001110111111011111010100001000111111101100111001000101100011011101111101101111011011101110011110111111110010100101000000110111110100000011000011101001011100001100010110000101011011010100100110111001001000100100101101000100101011000001011011000010000011000000101110101001100100001011110111101101100100111100011100100010100000011100100010100010010010110100100011100011100011000001111111001100111011100000111001110100111010010011011001100111000000111110100111100110100110010111111100000001001011110100101110100110111111000100110100111101111000110101111100101001100001011000000101000000011000111101010111111010100110101010001010001001110010010101100011011010110101001001111001011111001011110101101011010100110110111111110010000101100111000100010001110111111111101010110111110111100101010110011111100001110110000010010110011110111100100110000001111011011001110100000111001010111100000101100001001100101010001100101111110101110100100110101010010110100100110100011011101111100100001110011110110001100111110101000110101011101000001101110001110001100101011001010010101011011001100011100011111100100100101110010011011100101111000010111101001011110101000000100100100000001101111000011111101011111000101000000110010111101100010001111001111011000010100001000111011101010000011100101011010110001001111011000110100001110001110111010000000011100111100100101111010010001001110010101110011110101010010101001101101111100010011111110110101001011000010000011101111110010110100010010110010001001110100010100001011001011001111011101000000010000001101100001111100101010110000110010111010111010110000010101100011110000110110011011001111110010000100010110100010100010010000110000001110011101101000101000000011110010111010011100011110001101100110100001101011001101100010001011100010100010001001111110111111010000111000100101011011101001100011000110111101001001111011110100010011011110101101010001100001010111001111010011000000011111011100110000101000000011011111010111011000000000111000111101000101111001100110100010000000100001000011101110010001010100100101000010100001101101100001101100000000110100111100100110010111111100101101101111001000000100011111111010011110110100011100001011110011110010001100000011010001111011100010001101110011111000101110000111100001111101001011000000000110000001011001111010110011001100110010100110111111100001111100110110101001110000111100110100010110011101100001000100110101010100110111100001001000011011100101001010100001101001101010110010111011010011110000011101100001100011011101111110110110010101000001001100101100001111100101110001011100101000011011010011011111100110101111111000110100101000011001011001011010001011100110101101000001100011001000110000101101111111101011111110100101000010011100101010010010101011110001110111101001100110111101010110111111001000000110111100110110010111110011001101011000000001010001011011001111011100110000101001000101010111010011100011111000011001001001000101100100111011011000001100100110100111011101110001111101000101000101010101110011000011010100000100010110110010101111011111001001111111111110110011011010000111101100100100111011010111010100100001111000011010011101111101100011010000010110111110000011100110100010110011100111100001111101100101101110010010001011010101011101011000011110011010010011000011110111001111101011000010010101101101001011111011001101100011001111100001000010000000010000011011001011011001110001011110000010110011000110100000110110111001000100111000011101001011110111001111001011111011101010011111001010100110101100100010100011111000011100110111000010010110011010100100110101010110111110001111111111110111101111101011101001001001100100101100010001110011111101111110111011101001001001001011001010010010011011001111100101001010101011001011110100110001000111011100010100000100100111000101101000100000101101000110001100010110011110100001100001110001100111010011011000111111100011011001100100011110101001100100100011001111011001101010110010011100011101101101011100010010110101001111111111101001100011100100011101000001000101110110101010011100100000100100001101010011000010001000010100111101100100110111000110111010001011100001111011101110101101110000000100110001110010001100111110110010000110011010110000010011110001100100101101100010001000011011111100111111011110010000010001010110111001101011110101010010000011001111111110100000101101100111011101011010011001010101010100111101110110011110000000011111100011110111111001101011100111110101011001100110001100011100100010110010011010010100110010000110000010000100110001000010111110001011111100101010010000011010101111101100101110111100100101011010110000101001110100011001011100000110001000000011100011110100000001110000110010111100100111001001000100011010000011101000100101000001011100001010000011100110001101000101111100110110100011100101001110110101001111000101110000110111110000000000100011110100101101000000011011010001101001010001110000010100011011100110001011011100001000100010011101010011010110100011010101011110101110000101000000010110111111111010111100110001011110101010111101011001000100001001001101010110100010110101010001010100011010100001110001001001010000000010001000100100001011011010000101110001101111101011010100111101101101010001001101101000001011011011011101111111010111100111011011011101101001010111101010000101001110001111010101000010001001000101100000111011100000011011100001010110010100101010111011101101001100001111010111110001101111100000101001111110000001101111110110001010010011000101001100;
expected = 13560438;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);
#20;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd29;
noise_select = `BIG_N'b01011001111111110011101000101011010100011110001000001111101101110001001110111110011101111001011010110011101001000000011111101100000011101111010111100000011100100110111001111001011001000100001000001101001110010010111111110001111011101100010011101001001100010010100100110001111010111010011000100000110101001001100001000010000111001011001010101111110111010110010100010100101100110011011010010101011001010100100001101110101011011011101000100111010000111111000000011000100110001001001101011011100101010010101011000010111111111011100110100001100000001110010011010010111100011110100101110111011110011011101100110001011111011011111110101110101101011011101110001001010010001111111101111010001111110110110010101110001100111110100110110110000010111011101101000011111110011011111101001110110010011000001100111101110000110110101100001001000100101010000101010010101010100001110101100101100010000110000110101110111111110001110111110010000111000010101101000111101010010101001001100010001001110110010101011111000101000000011101011111010110101100011000001111010111011100101101111001000100000111100000110010100111111101100111010001100011100001011010110101111101010101100011001101000000111100100011111010001100110010001100110101111111001100101111010100011001110101100101101010101011001011011010011000000110011100010010111110011101100011110000111110001100100000100100110101110111001101101100000100000111110000010110101001001000001001101010100011110100100101100101011100110110010100101110000100101011000100001100001111001011101010001110100010110111000010000110010010110100000010110000110110100000111100110010111010110000110110101111110110101000000010100111010000100000011101010011000010101100111010111110110000111110011111101011101111011010010101011111101100100000011110110101011101011000111101010011110010000001110001010111011100100000110001101000011010010011110000010001111111010001001011010000111011110111100000111001101101001010100110101100101011001001100110010001001011101000111100100000111011001111011100100011101110000100111000100111101110110101111101011101010000001010110001101100101010000001001010101010111010100110111000111100010100101000100110001110001011011000000101011101100001101100111110110100001011001001100100010111101111011011001001010110010000000100111001011101010010111100110000111101101000100100111001011101111100010101101111110110111010100001001000111000001011010101111011011110011111100101100000011111010010110010001001001101110101100111000101011111011001101000111110110100001110011010100111010100000001110000101010011100001001101010101101001011110101011001010011110011000111000111110010110010010011111110011001001100100110010110110011100110001111000001001101011011011010100000101101001001101010001101100111111000001110011111011000010101101010000101011110101111110001011000010100110000001100000110000100011000110001000001000110001010011010010011100010000000011111110010101101101111101001101111001000001111010100000001001011100001010000110000001010011000101101001000101001010111100011010011100010001000110001100110000100001101111001100000101001000010110111100111111011100101101000100110101001101011011111110011110011110001010000001110011010101001011100000110111010110100000100000000101101101010110111110011010000101010110000101000010001101101000000110011011111101011100010101010010011001110011001011111110010000101100000011111100011001110111011110010010001100001111011111001111011101111010001010100111100010000100111010100101110010111000111000001111110010101011010011010000011101011101000000000101000110011111001010010110110000110000111101000101100000011100000000010101011101010110110111011101100001111101011111000000011010100000110110000000011101011100011111000110111111000001011000100001010101111111100100000001000110011001101111001111100001110110000101000010100000000000011101010010101001111010010111001101111010110011000001100110111011110101101100001001110011001101101000110010101101101111001100001111111101101000101110110110001010110101110000110111010111000000010111100001011001011000001010101111110010101000010100111111010111101011101001101100010001011111111010000111000000100000110000000000000000000111011001010010111111111001011100010111100110110100111000111101010011010110001001110111011100010110101010101111011001010001110111011011101000111101100101110110100111111111110011110010001110111001111000101101000111100010100101100000000111001110110110101011101111110001001000100100000001101001111101101001111010100110001001001100110101001111110100111110111000100000011010101001010100100100110010110010111011001101100111011110010011011010000111110010010101000001101010101110010101111101001011011101101010011101111100001110100011111110001011111000010011100110000101000100110110011011001110101011011100001010011000110011010110000101011000110100010010111101010001010111010111011011101000111111000111110000101110101000111111001111010001001110111110001111110101111111110110001010111010001010110111010001100000110100110111011111011000011101100001101001101001000111000010101101010010100011111101010010000000010001111001100010101111100000111111101011010101001100000111001101110110011100111001111111101110110111001011110101001001110110010000110000000010000100000100111011111101000000011011101000100100010111001010000000000011011001110000000000101000100000110011001001010110111111110111111110010001011110011110011111011101000101011010110110101010011001011100111101001101011000110011001111110010110000000111111100011100001110111010100000110001000111000001100001000010000101001101111111111100011001101010001101001101110100100010010111101101010101001100011110101000110010110111000100010100101110011000001000001011010101011001101101110011111100100011001011011010100011000100111001000110010011011110110111001100110101000111101110011011010000010101011101010001010000010000110010000001001110101011010010100111011101100100100011110101110001110100101000000001011010000111110010011111100000001111011101011101100100100011011010111111011001101000011001001010100110000110110101000011100111001110101111111001110111001101101110101011100011011000000001000001100011111111110110011000101101110111101100011110000000110010000101000000010000011000001010010110000010000010010010100100011011101001000001110000001100010110100110111110101101001010110000001000111101100101000001000001100100111100010011011011010111100011101011011101010010101000110010110100000001100011100101011000010010101101101110100010010111110001011000011110010011110000100010100010001111;
expected = 6472567;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);
#20;
row = 0;
plaintext = `PLAINTEXT_WIDTH'd30;
noise_select = `BIG_N'b00010011010000100011011011111011000110111111000000010011111111101010011001011101011100000001111101000111111000001000011101111000011010100111011111110000100001011000110111101110011011010110000111011011000011010000111110111110111001010011101100101111101010001100000011011111000001110110010101100000110111010000100001010011010010101000011100101101100111011110101000010001010011001010001001001100110110111000110011101101011001100010101110111100101100000111001011010011110101010110100100100101101010111101000001000001011101001100110111010110101100000011101110101101001101111100110110100111110000011111110000111011001010010100011100010111111000100010011001000100010100011011111100011101001010101011101000100011011001100111000011001110110001100011110001000110111000111110010011001110010001001111001010111000100111010000111000100110100110110111111010010011111101111101100011100110011111100110100110011111111101101011001001010101111000010011101011010110110001100000101010001101000101100011111011110111001001100000000001000000010010001010101010111111001010011010010100100101001010100000001100101000000011001110011010011001111010011010010000110000010101010101010001100001100001001110101000110001010000011001100111001101111011110101011001010000111000001000100101110100001100001011001101010100110011100110111100000011010010010100111011011101001011110101110010001001001010010000101110010100010111001111000110110100100111111000100110000101000011110100000100011110000111101000111111101001000011111011010101111011100111101000100001110110011001011001011010110011101101111010010011101001001001111100001111101101100001101101101100111111110010111001100011111000010011001000111000100000100000010000111011110001000110111000001010010000000111110101110010101111011001001101101111011011001011100010010101101101011100100111100011001111010011110111101111101010011000000000111010000010000001110000111100101001000111100011011111100010101001110001110101010100101110100010000011111100000000110001101110001111110100001001001100111100011101110001001101011010001000001000101011100011111111000101101010010101100011001010100110001000100000101001110011111110110000111000010111111101101111010000001011010011111100000010001101000100010010100000100000101000111011110101010011001111011111111010110111011101001011011111000010000001101111100101100110011001110111000101000001011110011111110000111011101111000101010011001000100110110001010111110001100100010110010101101111110111111100100000001100000101110110001001010111001011101010001010000100000110000011011101111111001000110010110110100011110101001010011111010010011101001100101001001010100100101111110100111101111100100101111101111010110111011110001011110011010011011110001010110011001101000000001101110101111010111001111101110000111111100011011111100000010000101001101110000000000001010011101111010010101010011011001000010110111000000010000111000011000110101100011001100001110100100000100110111110111010011111101111111111010101001100110100110011101000000101110111001011000001111101100101000111100011000000001101000100101111101111101101110111010110010000000110000100110011111100001101111011011101000001111001010111110110100000101010110000000000111101010110001011100010001101010010000000110111101000001010011010111010111000001111011111100010111110001001001010000011010011101101101111000010001001100000000000011011111100011010110011101000111010001110111001110100010001011001010110110001011111110100010101111100011111000000111010001110001111000111101011100110001110110011010111101001011000100110100110111011110111010000011001010100011000001011010110101010101000011100000101110011111101101111010001111100111001000010010001100111000000001001010111010111100010111110001100110011000000111111111110001001011000100101001110110101010100111111000011111010011110011001110010100001001001101100010010110111111011101000011111011000011100100000101100101111010001001001100001010000110000010111100011111110000101010100110110000111001000110010011110001110001000010101101100111001100011011000000011001000011100110110101011011101001110001010010011010000010011100101011100100100101110010111010110110100110111011001111100000010110001011001101010111100111011011001000010111100100001010100011100001001010111110111100011101011000011010100111110010101000101101111101101111000001010110110101001011001001000001100111001010101100111100011110010100011110110101011010000101101001110011110001001011010100000100101010100111111110111010111110101101000011100101001011111011000101000001001101110101111010011110111010001001011111000111010101100101110111101011000010110110101000011101111010001111111110010010010010100010110100011001011011010111010101100001000001100001011011100010101000010001001010000110000111011111110010010010000110101011001000110101010011010101110110110111001101111111101111101000111010010010010111000011110110000011100111011011001011000001000001111111101101100011101100000011101010100100001111110000111010111111111100010101110000000100110001100101011000100001001010010111111111111011110111010011001110000000010010011100100101011101000100100001100011010111001000000111000001100101000101000010101001110100110000011001111001010100101001110100001101011100000000110101001011010010110111011100001110111010010000000111111101101110011010101001001010000100000111101001110101001101101001000100011110111100110111100111110011100100010010011110101000100010011001001010010000010100100100110110001001000110011111000010000000101100111000101101101110010110000110011110010101010111010011100101110101111010011001010000001000111011001100111111011001101100111001110010111110001100011010111001111110010100001000010101111111001000000010011111000101110110011110110000001011011000111100011111011000111010000101010001110010101010010111110100011011110101101001001101100100100000101010100111111000101011000100100000100000100101010011011111110000000110111100011001101110011111011001000110110011001011000001111101101001110010100101101100001001001100011101110101010010010011010111010001100110110010001011111101010110101010111110010011100001111010000100100010010011110000001011001111110000101110011010110010000010000100010111111110101010000100000001010010011001010001010011111001100111100001001010011101011001100110010100010110110011000100001110110110100000110110111110000111011100110110110101110000110001101011111010011100100011011000101101110101100011101101011001111110011001000110011010001011010100110111110100011010110011110100110100111000100100000111110110101111;
expected = 14940967;
#20;
$display("Result = %d", ciphertext); assert(ciphertext == expected);

$finish;
end
endmodule
