../../6-sram/outputs/sky130_sram_1kbyte_1rw1r_32x256_8.lef