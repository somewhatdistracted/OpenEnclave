

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO top 
  PIN clk 
    ANTENNAPARTIALMETALAREA 0.4614 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.456 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.152 LAYER met4 ; 
    ANTENNAMAXAREACAR 9.15953 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 47.4913 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.114062 LAYER via4 ;
  END clk
  PIN rst_n 
    ANTENNAPARTIALMETALAREA 18.2562 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 97.832 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.6015 LAYER met4 ; 
    ANTENNAMAXAREACAR 77.0933 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 375.091 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.69315 LAYER via4 ;
  END rst_n
  PIN wb_clk_i 
    ANTENNAPARTIALMETALAREA 22.4322 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 120.104 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.477 LAYER met4 ; 
    ANTENNAMAXAREACAR 77.5688 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 404.384 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.05178 LAYER via4 ;
  END wb_clk_i
  PIN wb_rst_i 
    ANTENNAPARTIALMETALAREA 4.4604 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 23.784 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 8.3265 LAYER met4 ; 
    ANTENNAMAXAREACAR 21.9302 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 109.513 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.317271 LAYER via4 ;
  END wb_rst_i
  PIN wbs_stb_i 
    ANTENNAPARTIALMETALAREA 8.8044 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 46.952 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4 ; 
    ANTENNAMAXAREACAR 52.3097 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 278.307 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4 ;
  END wbs_stb_i
  PIN wbs_cyc_i 
    ANTENNAPARTIALMETALAREA 7.7064 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 41.096 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4 ; 
    ANTENNAMAXAREACAR 35.9594 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 190.17 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4 ;
  END wbs_cyc_i
  PIN wbs_we_i 
    ANTENNAPARTIALMETALAREA 0.855 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.496 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 59.1905 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 309.278 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_we_i
  PIN wbs_sel_i[3] 
  END wbs_sel_i[3]
  PIN wbs_sel_i[2] 
  END wbs_sel_i[2]
  PIN wbs_sel_i[1] 
  END wbs_sel_i[1]
  PIN wbs_sel_i[0] 
  END wbs_sel_i[0]
  PIN wbs_dat_i[31] 
    ANTENNAPARTIALMETALAREA 8.6214 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 45.976 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 73.4778 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 389.548 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_dat_i[31]
  PIN wbs_dat_i[30] 
    ANTENNAPARTIALMETALAREA 8.4384 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 45 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 79.5143 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 420.96 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_dat_i[30]
  PIN wbs_dat_i[29] 
    ANTENNAPARTIALMETALAREA 8.0724 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 43.048 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 72.7563 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 383.31 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_dat_i[29]
  PIN wbs_dat_i[28] 
    ANTENNAPARTIALMETALAREA 4.698 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 25.992 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 71.4944 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 376.802 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_dat_i[28]
  PIN wbs_dat_i[27] 
    ANTENNAPARTIALMETALAREA 8.6214 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 45.976 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 80.0071 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 421.659 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_dat_i[27]
  PIN wbs_dat_i[26] 
    ANTENNAPARTIALMETALAREA 7.1574 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 38.168 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 68.0734 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 354.278 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_dat_i[26]
  PIN wbs_dat_i[25] 
    ANTENNAPARTIALMETALAREA 8.0724 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 43.048 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 75.9881 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 400.183 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_dat_i[25]
  PIN wbs_dat_i[24] 
    ANTENNAPARTIALMETALAREA 8.6214 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 45.976 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 75.0246 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 397.278 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_dat_i[24]
  PIN wbs_dat_i[23] 
    ANTENNAPARTIALMETALAREA 8.175 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 44.536 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 91.3944 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 488.968 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_dat_i[23]
  PIN wbs_dat_i[22] 
    ANTENNAPARTIALMETALAREA 7.3984 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 35.328 LAYER met4 ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 5.872 LAYER met5 ;
    ANTENNAPARTIALMETALSIDEAREA 12.648 LAYER met5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met5 ; 
    ANTENNAMAXAREACAR 98.6127 LAYER met5 ;
    ANTENNAMAXSIDEAREACAR 346.69 LAYER met5 ;
  END wbs_dat_i[22]
  PIN wbs_dat_i[21] 
    ANTENNAPARTIALMETALAREA 7.3404 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 39.144 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 68.6032 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 360.77 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_dat_i[21]
  PIN wbs_dat_i[20] 
    ANTENNAPARTIALMETALAREA 8.6214 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 45.976 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 78.4738 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 413.992 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_dat_i[20]
  PIN wbs_dat_i[19] 
    ANTENNAPARTIALMETALAREA 5.2024 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 23.616 LAYER met4 ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 19.184 LAYER met5 ;
    ANTENNAPARTIALMETALSIDEAREA 40.296 LAYER met5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met5 ; 
    ANTENNAMAXAREACAR 190.813 LAYER met5 ;
    ANTENNAMAXSIDEAREACAR 491.349 LAYER met5 ;
  END wbs_dat_i[19]
  PIN wbs_dat_i[18] 
    ANTENNAPARTIALMETALAREA 8.6214 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 45.976 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 75.9183 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 401.214 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_dat_i[18]
  PIN wbs_dat_i[17] 
    ANTENNAPARTIALMETALAREA 0.2034 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.08 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 44.25 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 220.857 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_dat_i[17]
  PIN wbs_dat_i[16] 
    ANTENNAPARTIALMETALAREA 8.0724 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 43.048 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 78.3246 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 413.325 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_dat_i[16]
  PIN wbs_dat_i[15] 
    ANTENNAPARTIALMETALAREA 8.9874 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 47.928 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 83.4286 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 440.159 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_dat_i[15]
  PIN wbs_dat_i[14] 
    ANTENNAPARTIALMETALAREA 8.6214 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 45.976 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 79.7341 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 421.373 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_dat_i[14]
  PIN wbs_dat_i[13] 
    ANTENNAPARTIALMETALAREA 8.0724 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 43.048 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 76.3341 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 401.198 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_dat_i[13]
  PIN wbs_dat_i[12] 
    ANTENNAPARTIALMETALAREA 7.3404 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 39.144 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 68.7183 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 361.881 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_dat_i[12]
  PIN wbs_dat_i[11] 
    ANTENNAPARTIALMETALAREA 8.0724 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 43.048 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 72.8484 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 384.119 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_dat_i[11]
  PIN wbs_dat_i[10] 
    ANTENNAPARTIALMETALAREA 8.4384 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 45 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 76.6246 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 404.881 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_dat_i[10]
  PIN wbs_dat_i[9] 
    ANTENNAPARTIALMETALAREA 1.587 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.4 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 57.4849 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 299.984 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_dat_i[9]
  PIN wbs_dat_i[8] 
    ANTENNAPARTIALMETALAREA 2.709 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 15.384 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 66.1095 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 348.802 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_dat_i[8]
  PIN wbs_dat_i[7] 
    ANTENNAPARTIALMETALAREA 0.855 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.496 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 61.823 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 318.643 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_dat_i[7]
  PIN wbs_dat_i[6] 
    ANTENNAPARTIALMETALAREA 3.783 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 21.112 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 63.4754 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 333.556 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_dat_i[6]
  PIN wbs_dat_i[5] 
    ANTENNAPARTIALMETALAREA 1.953 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 11.352 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 63.5246 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 333.159 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_dat_i[5]
  PIN wbs_dat_i[4] 
    ANTENNAPARTIALMETALAREA 1.221 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.448 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 73.3357 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 380.825 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_dat_i[4]
  PIN wbs_dat_i[3] 
    ANTENNAPARTIALMETALAREA 4.332 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 24.04 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 64.546 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 342.722 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_dat_i[3]
  PIN wbs_dat_i[2] 
    ANTENNAPARTIALMETALAREA 3.234 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 18.184 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 63.5972 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 322.937 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_dat_i[2]
  PIN wbs_dat_i[1] 
    ANTENNAPARTIALMETALAREA 2.319 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 13.304 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 78.0643 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 406.071 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_dat_i[1]
  PIN wbs_dat_i[0] 
    ANTENNAPARTIALMETALAREA 2.685 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 15.256 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 106.781 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 543.976 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_dat_i[0]
  PIN wbs_adr_i[31] 
    ANTENNAPARTIALMETALAREA 1.587 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.4 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 70.9282 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 358.603 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_adr_i[31]
  PIN wbs_adr_i[30] 
    ANTENNAPARTIALMETALAREA 4.1424 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 22.088 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 129.885 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 668.77 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_adr_i[30]
  PIN wbs_adr_i[29] 
    ANTENNAPARTIALMETALAREA 9.2184 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 49.16 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4 ; 
    ANTENNAMAXAREACAR 90.6792 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 478.424 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4 ;
  END wbs_adr_i[29]
  PIN wbs_adr_i[28] 
    ANTENNAPARTIALMETALAREA 4.8264 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 25.736 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4 ; 
    ANTENNAMAXAREACAR 80.8723 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 423.79 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4 ;
  END wbs_adr_i[28]
  PIN wbs_adr_i[27] 
    ANTENNAPARTIALMETALAREA 6.0594 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 32.312 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 64.3516 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 334.087 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_adr_i[27]
  PIN wbs_adr_i[26] 
    ANTENNAPARTIALMETALAREA 8.4384 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 45 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 92.8361 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 490.96 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_adr_i[26]
  PIN wbs_adr_i[25] 
    ANTENNAPARTIALMETALAREA 8.2794 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 44.152 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 117.358 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 619.762 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_adr_i[25]
  PIN wbs_adr_i[24] 
    ANTENNAPARTIALMETALAREA 4.0464 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 21.576 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 76.1492 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 385.222 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_adr_i[24]
  PIN wbs_adr_i[23] 
    ANTENNAPARTIALMETALAREA 8.8044 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 46.952 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 80.3837 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 412.722 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_adr_i[23]
  PIN wbs_adr_i[22] 
    ANTENNAPARTIALMETALAREA 8.9874 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 47.928 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4 ; 
    ANTENNAMAXAREACAR 41.1624 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 215.115 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4 ;
  END wbs_adr_i[22]
  PIN wbs_adr_i[21] 
    ANTENNAPARTIALMETALAREA 8.6214 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 45.976 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ; 
    ANTENNAMAXAREACAR 113.275 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 593.508 LAYER met4 ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4 ;
  END wbs_adr_i[21]
  PIN wbs_adr_i[20] 
    ANTENNAPARTIALMETALAREA 7.7064 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 41.096 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4 ; 
    ANTENNAMAXAREACAR 54.0869 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 279.62 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4 ;
  END wbs_adr_i[20]
  PIN wbs_adr_i[19] 
    ANTENNAPARTIALMETALAREA 6.7914 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 36.216 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4 ; 
    ANTENNAMAXAREACAR 38.8085 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 203.632 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4 ;
  END wbs_adr_i[19]
  PIN wbs_adr_i[18] 
    ANTENNAPARTIALMETALAREA 6.7914 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 36.216 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4 ; 
    ANTENNAMAXAREACAR 41.087 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 211.248 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4 ;
  END wbs_adr_i[18]
  PIN wbs_adr_i[17] 
    ANTENNAPARTIALMETALAREA 6.7914 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 36.216 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4 ; 
    ANTENNAMAXAREACAR 43.3996 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 221.632 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4 ;
  END wbs_adr_i[17]
  PIN wbs_adr_i[16] 
    ANTENNAPARTIALMETALAREA 6.0594 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 32.312 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4 ; 
    ANTENNAMAXAREACAR 60.8457 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 318.525 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4 ;
  END wbs_adr_i[16]
  PIN wbs_adr_i[15] 
    ANTENNAPARTIALMETALAREA 6.7914 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 36.216 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4 ; 
    ANTENNAMAXAREACAR 42.4513 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 223.147 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4 ;
  END wbs_adr_i[15]
  PIN wbs_adr_i[14] 
    ANTENNAPARTIALMETALAREA 0.3864 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.056 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4 ; 
    ANTENNAMAXAREACAR 23.3447 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 112.424 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4 ;
  END wbs_adr_i[14]
  PIN wbs_adr_i[13] 
    ANTENNAPARTIALMETALAREA 5.3274 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 28.408 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4 ; 
    ANTENNAMAXAREACAR 44.5717 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 229.883 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4 ;
  END wbs_adr_i[13]
  PIN wbs_adr_i[12] 
    ANTENNAPARTIALMETALAREA 6.0594 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 32.312 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4 ; 
    ANTENNAMAXAREACAR 57.5002 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 300.683 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4 ;
  END wbs_adr_i[12]
  PIN wbs_adr_i[11] 
    ANTENNAPARTIALMETALAREA 4.7784 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 25.48 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4 ; 
    ANTENNAMAXAREACAR 91.1745 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 477.236 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4 ;
  END wbs_adr_i[11]
  PIN wbs_adr_i[10] 
    ANTENNAPARTIALMETALAREA 6.7914 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 36.216 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4 ; 
    ANTENNAMAXAREACAR 26.1736 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 138.196 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4 ;
  END wbs_adr_i[10]
  PIN wbs_adr_i[9] 
    ANTENNAPARTIALMETALAREA 8.6214 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 45.976 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4 ; 
    ANTENNAMAXAREACAR 17.4768 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 89.7498 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.315421 LAYER via4 ;
  END wbs_adr_i[9]
  PIN wbs_adr_i[8] 
    ANTENNAPARTIALMETALAREA 6.7914 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 36.216 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4 ; 
    ANTENNAMAXAREACAR 20.9349 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 104.734 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.315421 LAYER via4 ;
  END wbs_adr_i[8]
  PIN wbs_adr_i[7] 
    ANTENNAPARTIALMETALAREA 9.3534 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 49.88 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.825 LAYER met4 ; 
    ANTENNAMAXAREACAR 8.74914 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 43.4412 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.147674 LAYER via4 ;
  END wbs_adr_i[7]
  PIN wbs_adr_i[6] 
    ANTENNAPARTIALMETALAREA 18.2562 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 97.832 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5775 LAYER met4 ; 
    ANTENNAMAXAREACAR 60.3892 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 313.595 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.456964 LAYER via4 ;
  END wbs_adr_i[6]
  PIN wbs_adr_i[5] 
    ANTENNAPARTIALMETALAREA 4.2534 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 22.68 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5775 LAYER met4 ; 
    ANTENNAMAXAREACAR 79.849 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 406.622 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.367778 LAYER via4 ;
  END wbs_adr_i[5]
  PIN wbs_adr_i[4] 
    ANTENNAPARTIALMETALAREA 1.3014 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.936 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.4075 LAYER met4 ; 
    ANTENNAMAXAREACAR 24.4815 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 120.759 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.264515 LAYER via4 ;
  END wbs_adr_i[4]
  PIN wbs_adr_i[3] 
    ANTENNAPARTIALMETALAREA 4.4124 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 23.528 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5775 LAYER met4 ; 
    ANTENNAMAXAREACAR 36.7685 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 181.953 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.349299 LAYER via4 ;
  END wbs_adr_i[3]
  PIN wbs_adr_i[2] 
    ANTENNAPARTIALMETALAREA 6.0594 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 32.312 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5775 LAYER met4 ; 
    ANTENNAMAXAREACAR 18.4695 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 87.7004 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.25839 LAYER via4 ;
  END wbs_adr_i[2]
  PIN wbs_adr_i[1] 
    ANTENNAPARTIALMETALAREA 3.6804 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 19.624 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5775 LAYER met4 ; 
    ANTENNAMAXAREACAR 13.5082 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 64.4559 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.25839 LAYER via4 ;
  END wbs_adr_i[1]
  PIN wbs_adr_i[0] 
    ANTENNAPARTIALMETALAREA 6.0594 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 32.312 LAYER met4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.665 LAYER met4 ; 
    ANTENNAMAXAREACAR 12.2292 LAYER met4 ;
    ANTENNAMAXSIDEAREACAR 62.7519 LAYER met4 ;
    ANTENNAMAXCUTCAR 0.197594 LAYER via4 ;
  END wbs_adr_i[0]
  PIN wbs_ack_o 
    ANTENNADIFFAREA 0.429 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 0.2034 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.08 LAYER met4 ;
  END wbs_ack_o
  PIN wbs_dat_o[31] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 8.4384 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 45 LAYER met4 ;
  END wbs_dat_o[31]
  PIN wbs_dat_o[30] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 6.0594 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 32.312 LAYER met4 ;
  END wbs_dat_o[30]
  PIN wbs_dat_o[29] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 6.0594 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 32.312 LAYER met4 ;
  END wbs_dat_o[29]
  PIN wbs_dat_o[28] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 6.4254 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 34.264 LAYER met4 ;
  END wbs_dat_o[28]
  PIN wbs_dat_o[27] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 8.4384 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 45 LAYER met4 ;
  END wbs_dat_o[27]
  PIN wbs_dat_o[26] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 8.4384 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 45 LAYER met4 ;
  END wbs_dat_o[26]
  PIN wbs_dat_o[25] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 7.7064 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 41.096 LAYER met4 ;
  END wbs_dat_o[25]
  PIN wbs_dat_o[24] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 7.7064 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 41.096 LAYER met4 ;
  END wbs_dat_o[24]
  PIN wbs_dat_o[23] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 7.1574 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 38.168 LAYER met4 ;
  END wbs_dat_o[23]
  PIN wbs_dat_o[22] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 8.4384 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 45 LAYER met4 ;
  END wbs_dat_o[22]
  PIN wbs_dat_o[21] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 8.4384 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 45 LAYER met4 ;
  END wbs_dat_o[21]
  PIN wbs_dat_o[20] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 8.0724 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 43.048 LAYER met4 ;
  END wbs_dat_o[20]
  PIN wbs_dat_o[19] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 7.5234 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 40.12 LAYER met4 ;
  END wbs_dat_o[19]
  PIN wbs_dat_o[18] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 8.4384 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 45 LAYER met4 ;
  END wbs_dat_o[18]
  PIN wbs_dat_o[17] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 8.4384 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 45 LAYER met4 ;
  END wbs_dat_o[17]
  PIN wbs_dat_o[16] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 0.2034 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.08 LAYER met4 ;
  END wbs_dat_o[16]
  PIN wbs_dat_o[15] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 8.4384 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 45 LAYER met4 ;
  END wbs_dat_o[15]
  PIN wbs_dat_o[14] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 8.2554 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 44.024 LAYER met4 ;
  END wbs_dat_o[14]
  PIN wbs_dat_o[13] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 8.4384 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 45 LAYER met4 ;
  END wbs_dat_o[13]
  PIN wbs_dat_o[12] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 7.8894 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 42.072 LAYER met4 ;
  END wbs_dat_o[12]
  PIN wbs_dat_o[11] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 8.4384 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 45 LAYER met4 ;
  END wbs_dat_o[11]
  PIN wbs_dat_o[10] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 7.1574 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 38.168 LAYER met4 ;
  END wbs_dat_o[10]
  PIN wbs_dat_o[9] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 8.4384 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 45 LAYER met4 ;
  END wbs_dat_o[9]
  PIN wbs_dat_o[8] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 0.2034 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.08 LAYER met4 ;
  END wbs_dat_o[8]
  PIN wbs_dat_o[7] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 7.3404 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 39.144 LAYER met4 ;
  END wbs_dat_o[7]
  PIN wbs_dat_o[6] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 8.4384 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 45 LAYER met4 ;
  END wbs_dat_o[6]
  PIN wbs_dat_o[5] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 8.4384 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 45 LAYER met4 ;
  END wbs_dat_o[5]
  PIN wbs_dat_o[4] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 8.0724 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 43.048 LAYER met4 ;
  END wbs_dat_o[4]
  PIN wbs_dat_o[3] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 7.7064 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 41.096 LAYER met4 ;
  END wbs_dat_o[3]
  PIN wbs_dat_o[2] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 9.3534 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 49.88 LAYER met4 ;
  END wbs_dat_o[2]
  PIN wbs_dat_o[1] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 9.3534 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 49.88 LAYER met4 ;
  END wbs_dat_o[1]
  PIN wbs_dat_o[0] 
    ANTENNADIFFAREA 0.43675 LAYER met4 ; 
    ANTENNAPARTIALMETALAREA 10.8174 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 57.688 LAYER met4 ;
  END wbs_dat_o[0]
END top

END LIBRARY
