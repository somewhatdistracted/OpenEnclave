module sram
#(
    parameter DATA_WIDTH = 128,
    parameter ADDR_WIDTH = 10,
    parameter DEPTH = 1024
)
(
    input clk,
    input wen,
    input [ADDR_WIDTH - 1 : 0] wadr,
    input [DATA_WIDTH - 1 : 0] wdata,
    input ren,
    input [ADDR_WIDTH - 1 : 0] radr,
    output [DATA_WIDTH - 1 : 0] rdata
);

    genvar x, y;
    generate
        wire [DATA_WIDTH - 1 : 0] rdata_w [DEPTH/1024 - 1 : 0]; 
        reg  [ADDR_WIDTH - 1 : 0] radr_r;

        always @ (posedge clk) begin
            radr_r <= radr;
        end 

        for (x = 0; x < DATA_WIDTH/32; x = x + 1) begin: width_macro
            for (y = 0; y < DEPTH/256; y = y + 1) begin: depth_macro
                // note: Excerpted from EE272 Sram Wrapper:
                // note: The default behavioral model generated by OpenRAM has an arbitrary
                //       delay of 3ns. Since the SRAM data is only valid for half a cycle
                //       any delay < half a cycle will not affect the simulation result.
                //       Since we will try to push for a clock period of 5ns, we manually
                //       changed the delay number to 1ns (< 2.5ns) to prevent functional error.
                sky130_sram_1kbyte_1rw1r_32x256_8 sram (
                .clk0(clk),
                .csb0(~(wen && (wadr[ADDR_WIDTH - 1 : 8] == y))),
                .web0(~(wen && (wadr[ADDR_WIDTH - 1 : 8] == y))), // And wadr in range
                .wmask0(4'hF),
                .addr0(wadr[7:0]),
                .din0(wdata[32*(x+1)-1 : 32*x]),
                .dout0(),
                .clk1(clk),
                .csb1(~(ren && (radr[ADDR_WIDTH - 1 : 8] == y))), // And radr in range
                .addr1(radr[7:0]),
                .dout1(rdata_w[y][32*(x+1)-1 : 32*x])
                );
            end
        end

        assign rdata = rdata_w[radr_r[ADDR_WIDTH - 1 : 8]];

    endgenerate

endmodule
