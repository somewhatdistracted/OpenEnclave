`define PLAINTEXT_MODULUS 32
`define PLAINTEXT_WIDTH 5
`define DIMENSION 128
`define CIPHERTEXT_MODULUS 16777216
`define CIPHERTEXT_WIDTH 24
`define BIG_N 6425

module decrypt_tb;

    reg clk;
    reg rst_n;
    reg [`CIPHERTEXT_WIDTH-1:0] secret_key [`DIMENSION:0];
    reg signed [`CIPHERTEXT_WIDTH-1:0] cipher_text [`DIMENSION:0];
    reg [`CIPHERTEXT_WIDTH-1:0] skentry;
    reg signed [`CIPHERTEXT_WIDTH-1:0] ctentry;
    reg [`DIMENSION:0] row;
    wire [`PLAINTEXT_WIDTH-1:0] result;
    reg [`PLAINTEXT_WIDTH-1:0] expected;

    always #10 clk = ~clk;

    decrypt #(
        .PLAINTEXT_MODULUS(`PLAINTEXT_MODULUS),
        .PLAINTEXT_WIDTH(`PLAINTEXT_WIDTH),
        .CIPHERTEXT_MODULUS(`CIPHERTEXT_MODULUS),
        .CIPHERTEXT_WIDTH(`CIPHERTEXT_WIDTH),
        .DIMENSION(`DIMENSION),
        .BIG_N(`BIG_N)
    ) decrypt_inst (
        .clk(clk),
        .rst_n(rst_n),
        .secretkey_entry(skentry),
        .ciphertext_entry(ctentry),
        .row(row),
        .result(result)
    );

    initial begin
clk = 0;
secret_key[0] = `CIPHERTEXT_WIDTH'd1;
secret_key[1] = `CIPHERTEXT_WIDTH'd5885794;
secret_key[2] = `CIPHERTEXT_WIDTH'd16090509;
secret_key[3] = `CIPHERTEXT_WIDTH'd8465743;
secret_key[4] = `CIPHERTEXT_WIDTH'd3563952;
secret_key[5] = `CIPHERTEXT_WIDTH'd10598768;
secret_key[6] = `CIPHERTEXT_WIDTH'd4826292;
secret_key[7] = `CIPHERTEXT_WIDTH'd13890339;
secret_key[8] = `CIPHERTEXT_WIDTH'd12654815;
secret_key[9] = `CIPHERTEXT_WIDTH'd3883635;
secret_key[10] = `CIPHERTEXT_WIDTH'd10237667;
secret_key[11] = `CIPHERTEXT_WIDTH'd5137832;
secret_key[12] = `CIPHERTEXT_WIDTH'd5200327;
secret_key[13] = `CIPHERTEXT_WIDTH'd1854201;
secret_key[14] = `CIPHERTEXT_WIDTH'd2857528;
secret_key[15] = `CIPHERTEXT_WIDTH'd3725106;
secret_key[16] = `CIPHERTEXT_WIDTH'd4655940;
secret_key[17] = `CIPHERTEXT_WIDTH'd2440515;
secret_key[18] = `CIPHERTEXT_WIDTH'd4249943;
secret_key[19] = `CIPHERTEXT_WIDTH'd10463956;
secret_key[20] = `CIPHERTEXT_WIDTH'd16218474;
secret_key[21] = `CIPHERTEXT_WIDTH'd10751245;
secret_key[22] = `CIPHERTEXT_WIDTH'd12327440;
secret_key[23] = `CIPHERTEXT_WIDTH'd7590268;
secret_key[24] = `CIPHERTEXT_WIDTH'd5547881;
secret_key[25] = `CIPHERTEXT_WIDTH'd4441131;
secret_key[26] = `CIPHERTEXT_WIDTH'd11631794;
secret_key[27] = `CIPHERTEXT_WIDTH'd7064948;
secret_key[28] = `CIPHERTEXT_WIDTH'd15036162;
secret_key[29] = `CIPHERTEXT_WIDTH'd3042978;
secret_key[30] = `CIPHERTEXT_WIDTH'd10804389;
secret_key[31] = `CIPHERTEXT_WIDTH'd13353831;
secret_key[32] = `CIPHERTEXT_WIDTH'd16226060;
secret_key[33] = `CIPHERTEXT_WIDTH'd12016671;
secret_key[34] = `CIPHERTEXT_WIDTH'd4272433;
secret_key[35] = `CIPHERTEXT_WIDTH'd11537198;
secret_key[36] = `CIPHERTEXT_WIDTH'd1973740;
secret_key[37] = `CIPHERTEXT_WIDTH'd7704422;
secret_key[38] = `CIPHERTEXT_WIDTH'd7208992;
secret_key[39] = `CIPHERTEXT_WIDTH'd4352000;
secret_key[40] = `CIPHERTEXT_WIDTH'd9702637;
secret_key[41] = `CIPHERTEXT_WIDTH'd217513;
secret_key[42] = `CIPHERTEXT_WIDTH'd8781349;
secret_key[43] = `CIPHERTEXT_WIDTH'd15902478;
secret_key[44] = `CIPHERTEXT_WIDTH'd7866657;
secret_key[45] = `CIPHERTEXT_WIDTH'd7245081;
secret_key[46] = `CIPHERTEXT_WIDTH'd13983577;
secret_key[47] = `CIPHERTEXT_WIDTH'd9479851;
secret_key[48] = `CIPHERTEXT_WIDTH'd4854150;
secret_key[49] = `CIPHERTEXT_WIDTH'd26550;
secret_key[50] = `CIPHERTEXT_WIDTH'd11516466;
secret_key[51] = `CIPHERTEXT_WIDTH'd14424476;
secret_key[52] = `CIPHERTEXT_WIDTH'd14627784;
secret_key[53] = `CIPHERTEXT_WIDTH'd12024688;
secret_key[54] = `CIPHERTEXT_WIDTH'd1849459;
secret_key[55] = `CIPHERTEXT_WIDTH'd15616611;
secret_key[56] = `CIPHERTEXT_WIDTH'd8804613;
secret_key[57] = `CIPHERTEXT_WIDTH'd3322229;
secret_key[58] = `CIPHERTEXT_WIDTH'd15636975;
secret_key[59] = `CIPHERTEXT_WIDTH'd579739;
secret_key[60] = `CIPHERTEXT_WIDTH'd9477259;
secret_key[61] = `CIPHERTEXT_WIDTH'd4201176;
secret_key[62] = `CIPHERTEXT_WIDTH'd165969;
secret_key[63] = `CIPHERTEXT_WIDTH'd12433874;
secret_key[64] = `CIPHERTEXT_WIDTH'd8131838;
secret_key[65] = `CIPHERTEXT_WIDTH'd127642;
secret_key[66] = `CIPHERTEXT_WIDTH'd7855128;
secret_key[67] = `CIPHERTEXT_WIDTH'd169083;
secret_key[68] = `CIPHERTEXT_WIDTH'd1958998;
secret_key[69] = `CIPHERTEXT_WIDTH'd10233558;
secret_key[70] = `CIPHERTEXT_WIDTH'd4653543;
secret_key[71] = `CIPHERTEXT_WIDTH'd4971053;
secret_key[72] = `CIPHERTEXT_WIDTH'd12784878;
secret_key[73] = `CIPHERTEXT_WIDTH'd8984983;
secret_key[74] = `CIPHERTEXT_WIDTH'd204958;
secret_key[75] = `CIPHERTEXT_WIDTH'd5857954;
secret_key[76] = `CIPHERTEXT_WIDTH'd3350983;
secret_key[77] = `CIPHERTEXT_WIDTH'd10163002;
secret_key[78] = `CIPHERTEXT_WIDTH'd588198;
secret_key[79] = `CIPHERTEXT_WIDTH'd7793405;
secret_key[80] = `CIPHERTEXT_WIDTH'd8787718;
secret_key[81] = `CIPHERTEXT_WIDTH'd13319771;
secret_key[82] = `CIPHERTEXT_WIDTH'd2069151;
secret_key[83] = `CIPHERTEXT_WIDTH'd3914360;
secret_key[84] = `CIPHERTEXT_WIDTH'd3067235;
secret_key[85] = `CIPHERTEXT_WIDTH'd1514793;
secret_key[86] = `CIPHERTEXT_WIDTH'd14591785;
secret_key[87] = `CIPHERTEXT_WIDTH'd3870533;
secret_key[88] = `CIPHERTEXT_WIDTH'd14778772;
secret_key[89] = `CIPHERTEXT_WIDTH'd3419365;
secret_key[90] = `CIPHERTEXT_WIDTH'd4527201;
secret_key[91] = `CIPHERTEXT_WIDTH'd13192218;
secret_key[92] = `CIPHERTEXT_WIDTH'd7018618;
secret_key[93] = `CIPHERTEXT_WIDTH'd10427523;
secret_key[94] = `CIPHERTEXT_WIDTH'd7772661;
secret_key[95] = `CIPHERTEXT_WIDTH'd12333444;
secret_key[96] = `CIPHERTEXT_WIDTH'd2034072;
secret_key[97] = `CIPHERTEXT_WIDTH'd3049502;
secret_key[98] = `CIPHERTEXT_WIDTH'd8481617;
secret_key[99] = `CIPHERTEXT_WIDTH'd11087038;
secret_key[100] = `CIPHERTEXT_WIDTH'd3753111;
secret_key[101] = `CIPHERTEXT_WIDTH'd5401396;
secret_key[102] = `CIPHERTEXT_WIDTH'd12843149;
secret_key[103] = `CIPHERTEXT_WIDTH'd14219882;
secret_key[104] = `CIPHERTEXT_WIDTH'd12958011;
secret_key[105] = `CIPHERTEXT_WIDTH'd3488773;
secret_key[106] = `CIPHERTEXT_WIDTH'd9168153;
secret_key[107] = `CIPHERTEXT_WIDTH'd96590;
secret_key[108] = `CIPHERTEXT_WIDTH'd5700742;
secret_key[109] = `CIPHERTEXT_WIDTH'd4576872;
secret_key[110] = `CIPHERTEXT_WIDTH'd7178831;
secret_key[111] = `CIPHERTEXT_WIDTH'd4700175;
secret_key[112] = `CIPHERTEXT_WIDTH'd6675992;
secret_key[113] = `CIPHERTEXT_WIDTH'd302477;
secret_key[114] = `CIPHERTEXT_WIDTH'd16444875;
secret_key[115] = `CIPHERTEXT_WIDTH'd8846019;
secret_key[116] = `CIPHERTEXT_WIDTH'd16315629;
secret_key[117] = `CIPHERTEXT_WIDTH'd16116583;
secret_key[118] = `CIPHERTEXT_WIDTH'd7780318;
secret_key[119] = `CIPHERTEXT_WIDTH'd13729641;
secret_key[120] = `CIPHERTEXT_WIDTH'd337592;
secret_key[121] = `CIPHERTEXT_WIDTH'd9390982;
secret_key[122] = `CIPHERTEXT_WIDTH'd2445565;
secret_key[123] = `CIPHERTEXT_WIDTH'd14774167;
secret_key[124] = `CIPHERTEXT_WIDTH'd6855142;
secret_key[125] = `CIPHERTEXT_WIDTH'd12852194;
secret_key[126] = `CIPHERTEXT_WIDTH'd4064569;
secret_key[127] = `CIPHERTEXT_WIDTH'd3905551;
secret_key[128] = `CIPHERTEXT_WIDTH'd5758701;
expected = 0;
cipher_text[0] = `CIPHERTEXT_WIDTH'd2515365;
cipher_text[1] = `CIPHERTEXT_WIDTH'd12946660;
cipher_text[2] = `CIPHERTEXT_WIDTH'd619420;
cipher_text[3] = `CIPHERTEXT_WIDTH'd6930257;
cipher_text[4] = `CIPHERTEXT_WIDTH'd7740586;
cipher_text[5] = `CIPHERTEXT_WIDTH'd6499201;
cipher_text[6] = `CIPHERTEXT_WIDTH'd3595638;
cipher_text[7] = `CIPHERTEXT_WIDTH'd10803105;
cipher_text[8] = `CIPHERTEXT_WIDTH'd16550648;
cipher_text[9] = `CIPHERTEXT_WIDTH'd9854791;
cipher_text[10] = `CIPHERTEXT_WIDTH'd4996269;
cipher_text[11] = `CIPHERTEXT_WIDTH'd6827467;
cipher_text[12] = `CIPHERTEXT_WIDTH'd13039809;
cipher_text[13] = `CIPHERTEXT_WIDTH'd10891236;
cipher_text[14] = `CIPHERTEXT_WIDTH'd14299432;
cipher_text[15] = `CIPHERTEXT_WIDTH'd8610028;
cipher_text[16] = `CIPHERTEXT_WIDTH'd13869921;
cipher_text[17] = `CIPHERTEXT_WIDTH'd11502842;
cipher_text[18] = `CIPHERTEXT_WIDTH'd14663668;
cipher_text[19] = `CIPHERTEXT_WIDTH'd4972960;
cipher_text[20] = `CIPHERTEXT_WIDTH'd11431921;
cipher_text[21] = `CIPHERTEXT_WIDTH'd2572787;
cipher_text[22] = `CIPHERTEXT_WIDTH'd2792004;
cipher_text[23] = `CIPHERTEXT_WIDTH'd13262389;
cipher_text[24] = `CIPHERTEXT_WIDTH'd5844471;
cipher_text[25] = `CIPHERTEXT_WIDTH'd11282014;
cipher_text[26] = `CIPHERTEXT_WIDTH'd11743198;
cipher_text[27] = `CIPHERTEXT_WIDTH'd6895987;
cipher_text[28] = `CIPHERTEXT_WIDTH'd3622964;
cipher_text[29] = `CIPHERTEXT_WIDTH'd11157469;
cipher_text[30] = `CIPHERTEXT_WIDTH'd9752620;
cipher_text[31] = `CIPHERTEXT_WIDTH'd4224531;
cipher_text[32] = `CIPHERTEXT_WIDTH'd11335001;
cipher_text[33] = `CIPHERTEXT_WIDTH'd6885866;
cipher_text[34] = `CIPHERTEXT_WIDTH'd9216506;
cipher_text[35] = `CIPHERTEXT_WIDTH'd7542951;
cipher_text[36] = `CIPHERTEXT_WIDTH'd7290160;
cipher_text[37] = `CIPHERTEXT_WIDTH'd5526489;
cipher_text[38] = `CIPHERTEXT_WIDTH'd12669207;
cipher_text[39] = `CIPHERTEXT_WIDTH'd4882028;
cipher_text[40] = `CIPHERTEXT_WIDTH'd1323614;
cipher_text[41] = `CIPHERTEXT_WIDTH'd15833853;
cipher_text[42] = `CIPHERTEXT_WIDTH'd9538804;
cipher_text[43] = `CIPHERTEXT_WIDTH'd15088428;
cipher_text[44] = `CIPHERTEXT_WIDTH'd8490145;
cipher_text[45] = `CIPHERTEXT_WIDTH'd6653268;
cipher_text[46] = `CIPHERTEXT_WIDTH'd5810477;
cipher_text[47] = `CIPHERTEXT_WIDTH'd3938668;
cipher_text[48] = `CIPHERTEXT_WIDTH'd6837126;
cipher_text[49] = `CIPHERTEXT_WIDTH'd13750215;
cipher_text[50] = `CIPHERTEXT_WIDTH'd3557280;
cipher_text[51] = `CIPHERTEXT_WIDTH'd2512442;
cipher_text[52] = `CIPHERTEXT_WIDTH'd4024396;
cipher_text[53] = `CIPHERTEXT_WIDTH'd15029755;
cipher_text[54] = `CIPHERTEXT_WIDTH'd9157359;
cipher_text[55] = `CIPHERTEXT_WIDTH'd16438482;
cipher_text[56] = `CIPHERTEXT_WIDTH'd12563241;
cipher_text[57] = `CIPHERTEXT_WIDTH'd712790;
cipher_text[58] = `CIPHERTEXT_WIDTH'd3175264;
cipher_text[59] = `CIPHERTEXT_WIDTH'd1546323;
cipher_text[60] = `CIPHERTEXT_WIDTH'd11889568;
cipher_text[61] = `CIPHERTEXT_WIDTH'd12558406;
cipher_text[62] = `CIPHERTEXT_WIDTH'd11744915;
cipher_text[63] = `CIPHERTEXT_WIDTH'd2471142;
cipher_text[64] = `CIPHERTEXT_WIDTH'd405052;
cipher_text[65] = `CIPHERTEXT_WIDTH'd7667783;
cipher_text[66] = `CIPHERTEXT_WIDTH'd15084741;
cipher_text[67] = `CIPHERTEXT_WIDTH'd12575515;
cipher_text[68] = `CIPHERTEXT_WIDTH'd11064288;
cipher_text[69] = `CIPHERTEXT_WIDTH'd11205166;
cipher_text[70] = `CIPHERTEXT_WIDTH'd14117546;
cipher_text[71] = `CIPHERTEXT_WIDTH'd4433811;
cipher_text[72] = `CIPHERTEXT_WIDTH'd9094475;
cipher_text[73] = `CIPHERTEXT_WIDTH'd9149370;
cipher_text[74] = `CIPHERTEXT_WIDTH'd14118558;
cipher_text[75] = `CIPHERTEXT_WIDTH'd13152199;
cipher_text[76] = `CIPHERTEXT_WIDTH'd11820690;
cipher_text[77] = `CIPHERTEXT_WIDTH'd12316132;
cipher_text[78] = `CIPHERTEXT_WIDTH'd15246235;
cipher_text[79] = `CIPHERTEXT_WIDTH'd10094201;
cipher_text[80] = `CIPHERTEXT_WIDTH'd5203532;
cipher_text[81] = `CIPHERTEXT_WIDTH'd14955225;
cipher_text[82] = `CIPHERTEXT_WIDTH'd15369000;
cipher_text[83] = `CIPHERTEXT_WIDTH'd14662445;
cipher_text[84] = `CIPHERTEXT_WIDTH'd10737445;
cipher_text[85] = `CIPHERTEXT_WIDTH'd11437031;
cipher_text[86] = `CIPHERTEXT_WIDTH'd14399727;
cipher_text[87] = `CIPHERTEXT_WIDTH'd7369027;
cipher_text[88] = `CIPHERTEXT_WIDTH'd9175448;
cipher_text[89] = `CIPHERTEXT_WIDTH'd6984920;
cipher_text[90] = `CIPHERTEXT_WIDTH'd5030723;
cipher_text[91] = `CIPHERTEXT_WIDTH'd706535;
cipher_text[92] = `CIPHERTEXT_WIDTH'd2035497;
cipher_text[93] = `CIPHERTEXT_WIDTH'd9418696;
cipher_text[94] = `CIPHERTEXT_WIDTH'd11098975;
cipher_text[95] = `CIPHERTEXT_WIDTH'd512955;
cipher_text[96] = `CIPHERTEXT_WIDTH'd2573606;
cipher_text[97] = `CIPHERTEXT_WIDTH'd9357477;
cipher_text[98] = `CIPHERTEXT_WIDTH'd3659425;
cipher_text[99] = `CIPHERTEXT_WIDTH'd13226920;
cipher_text[100] = `CIPHERTEXT_WIDTH'd7613942;
cipher_text[101] = `CIPHERTEXT_WIDTH'd7929203;
cipher_text[102] = `CIPHERTEXT_WIDTH'd9044662;
cipher_text[103] = `CIPHERTEXT_WIDTH'd15144479;
cipher_text[104] = `CIPHERTEXT_WIDTH'd317630;
cipher_text[105] = `CIPHERTEXT_WIDTH'd6003380;
cipher_text[106] = `CIPHERTEXT_WIDTH'd10020100;
cipher_text[107] = `CIPHERTEXT_WIDTH'd13795903;
cipher_text[108] = `CIPHERTEXT_WIDTH'd7463190;
cipher_text[109] = `CIPHERTEXT_WIDTH'd6806914;
cipher_text[110] = `CIPHERTEXT_WIDTH'd8898519;
cipher_text[111] = `CIPHERTEXT_WIDTH'd1677870;
cipher_text[112] = `CIPHERTEXT_WIDTH'd4442947;
cipher_text[113] = `CIPHERTEXT_WIDTH'd14641771;
cipher_text[114] = `CIPHERTEXT_WIDTH'd11039089;
cipher_text[115] = `CIPHERTEXT_WIDTH'd10729955;
cipher_text[116] = `CIPHERTEXT_WIDTH'd16182329;
cipher_text[117] = `CIPHERTEXT_WIDTH'd4822185;
cipher_text[118] = `CIPHERTEXT_WIDTH'd12839769;
cipher_text[119] = `CIPHERTEXT_WIDTH'd9076877;
cipher_text[120] = `CIPHERTEXT_WIDTH'd12029828;
cipher_text[121] = `CIPHERTEXT_WIDTH'd6597177;
cipher_text[122] = `CIPHERTEXT_WIDTH'd3125067;
cipher_text[123] = `CIPHERTEXT_WIDTH'd2924545;
cipher_text[124] = `CIPHERTEXT_WIDTH'd1120678;
cipher_text[125] = `CIPHERTEXT_WIDTH'd7077870;
cipher_text[126] = `CIPHERTEXT_WIDTH'd5530095;
cipher_text[127] = `CIPHERTEXT_WIDTH'd16488999;
cipher_text[128] = `CIPHERTEXT_WIDTH'd780360;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 1;
cipher_text[0] = `CIPHERTEXT_WIDTH'd12090373;
cipher_text[1] = `CIPHERTEXT_WIDTH'd16494165;
cipher_text[2] = `CIPHERTEXT_WIDTH'd15906125;
cipher_text[3] = `CIPHERTEXT_WIDTH'd11789969;
cipher_text[4] = `CIPHERTEXT_WIDTH'd179039;
cipher_text[5] = `CIPHERTEXT_WIDTH'd7383896;
cipher_text[6] = `CIPHERTEXT_WIDTH'd4100808;
cipher_text[7] = `CIPHERTEXT_WIDTH'd2620256;
cipher_text[8] = `CIPHERTEXT_WIDTH'd9767969;
cipher_text[9] = `CIPHERTEXT_WIDTH'd7884427;
cipher_text[10] = `CIPHERTEXT_WIDTH'd2175681;
cipher_text[11] = `CIPHERTEXT_WIDTH'd5711006;
cipher_text[12] = `CIPHERTEXT_WIDTH'd1690208;
cipher_text[13] = `CIPHERTEXT_WIDTH'd13275451;
cipher_text[14] = `CIPHERTEXT_WIDTH'd3319153;
cipher_text[15] = `CIPHERTEXT_WIDTH'd9484682;
cipher_text[16] = `CIPHERTEXT_WIDTH'd8144238;
cipher_text[17] = `CIPHERTEXT_WIDTH'd3678704;
cipher_text[18] = `CIPHERTEXT_WIDTH'd13625423;
cipher_text[19] = `CIPHERTEXT_WIDTH'd7342475;
cipher_text[20] = `CIPHERTEXT_WIDTH'd3841372;
cipher_text[21] = `CIPHERTEXT_WIDTH'd11827765;
cipher_text[22] = `CIPHERTEXT_WIDTH'd3707542;
cipher_text[23] = `CIPHERTEXT_WIDTH'd1225080;
cipher_text[24] = `CIPHERTEXT_WIDTH'd3319490;
cipher_text[25] = `CIPHERTEXT_WIDTH'd15323583;
cipher_text[26] = `CIPHERTEXT_WIDTH'd15020211;
cipher_text[27] = `CIPHERTEXT_WIDTH'd1904186;
cipher_text[28] = `CIPHERTEXT_WIDTH'd7858187;
cipher_text[29] = `CIPHERTEXT_WIDTH'd8431397;
cipher_text[30] = `CIPHERTEXT_WIDTH'd10149400;
cipher_text[31] = `CIPHERTEXT_WIDTH'd14549943;
cipher_text[32] = `CIPHERTEXT_WIDTH'd6694393;
cipher_text[33] = `CIPHERTEXT_WIDTH'd11155737;
cipher_text[34] = `CIPHERTEXT_WIDTH'd8152155;
cipher_text[35] = `CIPHERTEXT_WIDTH'd2007768;
cipher_text[36] = `CIPHERTEXT_WIDTH'd2133006;
cipher_text[37] = `CIPHERTEXT_WIDTH'd15215976;
cipher_text[38] = `CIPHERTEXT_WIDTH'd9954100;
cipher_text[39] = `CIPHERTEXT_WIDTH'd14343079;
cipher_text[40] = `CIPHERTEXT_WIDTH'd3548264;
cipher_text[41] = `CIPHERTEXT_WIDTH'd12895385;
cipher_text[42] = `CIPHERTEXT_WIDTH'd3691792;
cipher_text[43] = `CIPHERTEXT_WIDTH'd7890835;
cipher_text[44] = `CIPHERTEXT_WIDTH'd5501216;
cipher_text[45] = `CIPHERTEXT_WIDTH'd2865321;
cipher_text[46] = `CIPHERTEXT_WIDTH'd15797863;
cipher_text[47] = `CIPHERTEXT_WIDTH'd738084;
cipher_text[48] = `CIPHERTEXT_WIDTH'd3544205;
cipher_text[49] = `CIPHERTEXT_WIDTH'd6588797;
cipher_text[50] = `CIPHERTEXT_WIDTH'd10920584;
cipher_text[51] = `CIPHERTEXT_WIDTH'd566217;
cipher_text[52] = `CIPHERTEXT_WIDTH'd2748523;
cipher_text[53] = `CIPHERTEXT_WIDTH'd4261301;
cipher_text[54] = `CIPHERTEXT_WIDTH'd10488060;
cipher_text[55] = `CIPHERTEXT_WIDTH'd10789677;
cipher_text[56] = `CIPHERTEXT_WIDTH'd3096102;
cipher_text[57] = `CIPHERTEXT_WIDTH'd13885368;
cipher_text[58] = `CIPHERTEXT_WIDTH'd511181;
cipher_text[59] = `CIPHERTEXT_WIDTH'd14557936;
cipher_text[60] = `CIPHERTEXT_WIDTH'd12408187;
cipher_text[61] = `CIPHERTEXT_WIDTH'd3248362;
cipher_text[62] = `CIPHERTEXT_WIDTH'd3198993;
cipher_text[63] = `CIPHERTEXT_WIDTH'd9117608;
cipher_text[64] = `CIPHERTEXT_WIDTH'd15937148;
cipher_text[65] = `CIPHERTEXT_WIDTH'd13877157;
cipher_text[66] = `CIPHERTEXT_WIDTH'd14890364;
cipher_text[67] = `CIPHERTEXT_WIDTH'd15344719;
cipher_text[68] = `CIPHERTEXT_WIDTH'd1606859;
cipher_text[69] = `CIPHERTEXT_WIDTH'd11924253;
cipher_text[70] = `CIPHERTEXT_WIDTH'd15502703;
cipher_text[71] = `CIPHERTEXT_WIDTH'd6650262;
cipher_text[72] = `CIPHERTEXT_WIDTH'd10002867;
cipher_text[73] = `CIPHERTEXT_WIDTH'd14046033;
cipher_text[74] = `CIPHERTEXT_WIDTH'd10803045;
cipher_text[75] = `CIPHERTEXT_WIDTH'd4490020;
cipher_text[76] = `CIPHERTEXT_WIDTH'd537556;
cipher_text[77] = `CIPHERTEXT_WIDTH'd10018613;
cipher_text[78] = `CIPHERTEXT_WIDTH'd12270789;
cipher_text[79] = `CIPHERTEXT_WIDTH'd8919451;
cipher_text[80] = `CIPHERTEXT_WIDTH'd1947645;
cipher_text[81] = `CIPHERTEXT_WIDTH'd14615474;
cipher_text[82] = `CIPHERTEXT_WIDTH'd15377070;
cipher_text[83] = `CIPHERTEXT_WIDTH'd13250461;
cipher_text[84] = `CIPHERTEXT_WIDTH'd4142387;
cipher_text[85] = `CIPHERTEXT_WIDTH'd5910363;
cipher_text[86] = `CIPHERTEXT_WIDTH'd1544816;
cipher_text[87] = `CIPHERTEXT_WIDTH'd157341;
cipher_text[88] = `CIPHERTEXT_WIDTH'd11095117;
cipher_text[89] = `CIPHERTEXT_WIDTH'd12516486;
cipher_text[90] = `CIPHERTEXT_WIDTH'd11657941;
cipher_text[91] = `CIPHERTEXT_WIDTH'd2954944;
cipher_text[92] = `CIPHERTEXT_WIDTH'd9875979;
cipher_text[93] = `CIPHERTEXT_WIDTH'd433685;
cipher_text[94] = `CIPHERTEXT_WIDTH'd1344278;
cipher_text[95] = `CIPHERTEXT_WIDTH'd7147902;
cipher_text[96] = `CIPHERTEXT_WIDTH'd2592472;
cipher_text[97] = `CIPHERTEXT_WIDTH'd3646862;
cipher_text[98] = `CIPHERTEXT_WIDTH'd13250586;
cipher_text[99] = `CIPHERTEXT_WIDTH'd15124708;
cipher_text[100] = `CIPHERTEXT_WIDTH'd2983363;
cipher_text[101] = `CIPHERTEXT_WIDTH'd8265825;
cipher_text[102] = `CIPHERTEXT_WIDTH'd14295634;
cipher_text[103] = `CIPHERTEXT_WIDTH'd4077293;
cipher_text[104] = `CIPHERTEXT_WIDTH'd4162531;
cipher_text[105] = `CIPHERTEXT_WIDTH'd6519307;
cipher_text[106] = `CIPHERTEXT_WIDTH'd5565491;
cipher_text[107] = `CIPHERTEXT_WIDTH'd8876111;
cipher_text[108] = `CIPHERTEXT_WIDTH'd5446375;
cipher_text[109] = `CIPHERTEXT_WIDTH'd773784;
cipher_text[110] = `CIPHERTEXT_WIDTH'd10325768;
cipher_text[111] = `CIPHERTEXT_WIDTH'd6979381;
cipher_text[112] = `CIPHERTEXT_WIDTH'd7597391;
cipher_text[113] = `CIPHERTEXT_WIDTH'd4964138;
cipher_text[114] = `CIPHERTEXT_WIDTH'd8004453;
cipher_text[115] = `CIPHERTEXT_WIDTH'd10218266;
cipher_text[116] = `CIPHERTEXT_WIDTH'd7080607;
cipher_text[117] = `CIPHERTEXT_WIDTH'd2290874;
cipher_text[118] = `CIPHERTEXT_WIDTH'd9949261;
cipher_text[119] = `CIPHERTEXT_WIDTH'd12792508;
cipher_text[120] = `CIPHERTEXT_WIDTH'd8425724;
cipher_text[121] = `CIPHERTEXT_WIDTH'd3488434;
cipher_text[122] = `CIPHERTEXT_WIDTH'd10894573;
cipher_text[123] = `CIPHERTEXT_WIDTH'd6103820;
cipher_text[124] = `CIPHERTEXT_WIDTH'd12595105;
cipher_text[125] = `CIPHERTEXT_WIDTH'd14747498;
cipher_text[126] = `CIPHERTEXT_WIDTH'd635064;
cipher_text[127] = `CIPHERTEXT_WIDTH'd4723121;
cipher_text[128] = `CIPHERTEXT_WIDTH'd12098215;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 2;
cipher_text[0] = `CIPHERTEXT_WIDTH'd5141654;
cipher_text[1] = `CIPHERTEXT_WIDTH'd1546919;
cipher_text[2] = `CIPHERTEXT_WIDTH'd13268581;
cipher_text[3] = `CIPHERTEXT_WIDTH'd12613103;
cipher_text[4] = `CIPHERTEXT_WIDTH'd2673397;
cipher_text[5] = `CIPHERTEXT_WIDTH'd7245296;
cipher_text[6] = `CIPHERTEXT_WIDTH'd8283970;
cipher_text[7] = `CIPHERTEXT_WIDTH'd1498532;
cipher_text[8] = `CIPHERTEXT_WIDTH'd11407382;
cipher_text[9] = `CIPHERTEXT_WIDTH'd12709810;
cipher_text[10] = `CIPHERTEXT_WIDTH'd8561621;
cipher_text[11] = `CIPHERTEXT_WIDTH'd11549847;
cipher_text[12] = `CIPHERTEXT_WIDTH'd9018222;
cipher_text[13] = `CIPHERTEXT_WIDTH'd7912637;
cipher_text[14] = `CIPHERTEXT_WIDTH'd11452504;
cipher_text[15] = `CIPHERTEXT_WIDTH'd6429613;
cipher_text[16] = `CIPHERTEXT_WIDTH'd5805055;
cipher_text[17] = `CIPHERTEXT_WIDTH'd4545542;
cipher_text[18] = `CIPHERTEXT_WIDTH'd9066868;
cipher_text[19] = `CIPHERTEXT_WIDTH'd15380047;
cipher_text[20] = `CIPHERTEXT_WIDTH'd12186118;
cipher_text[21] = `CIPHERTEXT_WIDTH'd7557506;
cipher_text[22] = `CIPHERTEXT_WIDTH'd11563577;
cipher_text[23] = `CIPHERTEXT_WIDTH'd9084535;
cipher_text[24] = `CIPHERTEXT_WIDTH'd11149979;
cipher_text[25] = `CIPHERTEXT_WIDTH'd14615961;
cipher_text[26] = `CIPHERTEXT_WIDTH'd10258628;
cipher_text[27] = `CIPHERTEXT_WIDTH'd6625008;
cipher_text[28] = `CIPHERTEXT_WIDTH'd4395322;
cipher_text[29] = `CIPHERTEXT_WIDTH'd8821975;
cipher_text[30] = `CIPHERTEXT_WIDTH'd1800273;
cipher_text[31] = `CIPHERTEXT_WIDTH'd2102294;
cipher_text[32] = `CIPHERTEXT_WIDTH'd13124558;
cipher_text[33] = `CIPHERTEXT_WIDTH'd14131634;
cipher_text[34] = `CIPHERTEXT_WIDTH'd5236881;
cipher_text[35] = `CIPHERTEXT_WIDTH'd15019501;
cipher_text[36] = `CIPHERTEXT_WIDTH'd16751384;
cipher_text[37] = `CIPHERTEXT_WIDTH'd1144394;
cipher_text[38] = `CIPHERTEXT_WIDTH'd8167656;
cipher_text[39] = `CIPHERTEXT_WIDTH'd12123468;
cipher_text[40] = `CIPHERTEXT_WIDTH'd16084822;
cipher_text[41] = `CIPHERTEXT_WIDTH'd16303910;
cipher_text[42] = `CIPHERTEXT_WIDTH'd6644124;
cipher_text[43] = `CIPHERTEXT_WIDTH'd4749471;
cipher_text[44] = `CIPHERTEXT_WIDTH'd7719921;
cipher_text[45] = `CIPHERTEXT_WIDTH'd1400428;
cipher_text[46] = `CIPHERTEXT_WIDTH'd9832406;
cipher_text[47] = `CIPHERTEXT_WIDTH'd10828561;
cipher_text[48] = `CIPHERTEXT_WIDTH'd14951221;
cipher_text[49] = `CIPHERTEXT_WIDTH'd12684192;
cipher_text[50] = `CIPHERTEXT_WIDTH'd777102;
cipher_text[51] = `CIPHERTEXT_WIDTH'd5836581;
cipher_text[52] = `CIPHERTEXT_WIDTH'd655937;
cipher_text[53] = `CIPHERTEXT_WIDTH'd16265066;
cipher_text[54] = `CIPHERTEXT_WIDTH'd13068396;
cipher_text[55] = `CIPHERTEXT_WIDTH'd14757605;
cipher_text[56] = `CIPHERTEXT_WIDTH'd3615872;
cipher_text[57] = `CIPHERTEXT_WIDTH'd12278874;
cipher_text[58] = `CIPHERTEXT_WIDTH'd10572955;
cipher_text[59] = `CIPHERTEXT_WIDTH'd10525329;
cipher_text[60] = `CIPHERTEXT_WIDTH'd2588036;
cipher_text[61] = `CIPHERTEXT_WIDTH'd12407986;
cipher_text[62] = `CIPHERTEXT_WIDTH'd15299013;
cipher_text[63] = `CIPHERTEXT_WIDTH'd11525815;
cipher_text[64] = `CIPHERTEXT_WIDTH'd12688671;
cipher_text[65] = `CIPHERTEXT_WIDTH'd6685635;
cipher_text[66] = `CIPHERTEXT_WIDTH'd8136707;
cipher_text[67] = `CIPHERTEXT_WIDTH'd4980447;
cipher_text[68] = `CIPHERTEXT_WIDTH'd12463669;
cipher_text[69] = `CIPHERTEXT_WIDTH'd10360526;
cipher_text[70] = `CIPHERTEXT_WIDTH'd9434987;
cipher_text[71] = `CIPHERTEXT_WIDTH'd10780240;
cipher_text[72] = `CIPHERTEXT_WIDTH'd7310408;
cipher_text[73] = `CIPHERTEXT_WIDTH'd14585024;
cipher_text[74] = `CIPHERTEXT_WIDTH'd14394073;
cipher_text[75] = `CIPHERTEXT_WIDTH'd9982414;
cipher_text[76] = `CIPHERTEXT_WIDTH'd3807764;
cipher_text[77] = `CIPHERTEXT_WIDTH'd200448;
cipher_text[78] = `CIPHERTEXT_WIDTH'd9341287;
cipher_text[79] = `CIPHERTEXT_WIDTH'd12210471;
cipher_text[80] = `CIPHERTEXT_WIDTH'd5067395;
cipher_text[81] = `CIPHERTEXT_WIDTH'd10514866;
cipher_text[82] = `CIPHERTEXT_WIDTH'd10853174;
cipher_text[83] = `CIPHERTEXT_WIDTH'd1909441;
cipher_text[84] = `CIPHERTEXT_WIDTH'd11457082;
cipher_text[85] = `CIPHERTEXT_WIDTH'd16120671;
cipher_text[86] = `CIPHERTEXT_WIDTH'd7703570;
cipher_text[87] = `CIPHERTEXT_WIDTH'd15846914;
cipher_text[88] = `CIPHERTEXT_WIDTH'd8968853;
cipher_text[89] = `CIPHERTEXT_WIDTH'd6188020;
cipher_text[90] = `CIPHERTEXT_WIDTH'd13206550;
cipher_text[91] = `CIPHERTEXT_WIDTH'd3147935;
cipher_text[92] = `CIPHERTEXT_WIDTH'd10170113;
cipher_text[93] = `CIPHERTEXT_WIDTH'd2685441;
cipher_text[94] = `CIPHERTEXT_WIDTH'd11309119;
cipher_text[95] = `CIPHERTEXT_WIDTH'd11976110;
cipher_text[96] = `CIPHERTEXT_WIDTH'd2204102;
cipher_text[97] = `CIPHERTEXT_WIDTH'd5030263;
cipher_text[98] = `CIPHERTEXT_WIDTH'd8220696;
cipher_text[99] = `CIPHERTEXT_WIDTH'd13457235;
cipher_text[100] = `CIPHERTEXT_WIDTH'd8391344;
cipher_text[101] = `CIPHERTEXT_WIDTH'd5416279;
cipher_text[102] = `CIPHERTEXT_WIDTH'd7644744;
cipher_text[103] = `CIPHERTEXT_WIDTH'd10323080;
cipher_text[104] = `CIPHERTEXT_WIDTH'd16426300;
cipher_text[105] = `CIPHERTEXT_WIDTH'd10568413;
cipher_text[106] = `CIPHERTEXT_WIDTH'd14369433;
cipher_text[107] = `CIPHERTEXT_WIDTH'd7735844;
cipher_text[108] = `CIPHERTEXT_WIDTH'd6530292;
cipher_text[109] = `CIPHERTEXT_WIDTH'd7848133;
cipher_text[110] = `CIPHERTEXT_WIDTH'd1003400;
cipher_text[111] = `CIPHERTEXT_WIDTH'd13398103;
cipher_text[112] = `CIPHERTEXT_WIDTH'd9156902;
cipher_text[113] = `CIPHERTEXT_WIDTH'd9186954;
cipher_text[114] = `CIPHERTEXT_WIDTH'd7606219;
cipher_text[115] = `CIPHERTEXT_WIDTH'd12866869;
cipher_text[116] = `CIPHERTEXT_WIDTH'd3489280;
cipher_text[117] = `CIPHERTEXT_WIDTH'd9219176;
cipher_text[118] = `CIPHERTEXT_WIDTH'd3242290;
cipher_text[119] = `CIPHERTEXT_WIDTH'd1579836;
cipher_text[120] = `CIPHERTEXT_WIDTH'd12401083;
cipher_text[121] = `CIPHERTEXT_WIDTH'd1623833;
cipher_text[122] = `CIPHERTEXT_WIDTH'd4426329;
cipher_text[123] = `CIPHERTEXT_WIDTH'd15417944;
cipher_text[124] = `CIPHERTEXT_WIDTH'd6770388;
cipher_text[125] = `CIPHERTEXT_WIDTH'd16354287;
cipher_text[126] = `CIPHERTEXT_WIDTH'd5344837;
cipher_text[127] = `CIPHERTEXT_WIDTH'd5793057;
cipher_text[128] = `CIPHERTEXT_WIDTH'd16609578;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 3;
cipher_text[0] = `CIPHERTEXT_WIDTH'd16106645;
cipher_text[1] = `CIPHERTEXT_WIDTH'd13682922;
cipher_text[2] = `CIPHERTEXT_WIDTH'd12424817;
cipher_text[3] = `CIPHERTEXT_WIDTH'd15670222;
cipher_text[4] = `CIPHERTEXT_WIDTH'd5221874;
cipher_text[5] = `CIPHERTEXT_WIDTH'd13767844;
cipher_text[6] = `CIPHERTEXT_WIDTH'd16136284;
cipher_text[7] = `CIPHERTEXT_WIDTH'd7266118;
cipher_text[8] = `CIPHERTEXT_WIDTH'd2980975;
cipher_text[9] = `CIPHERTEXT_WIDTH'd15108100;
cipher_text[10] = `CIPHERTEXT_WIDTH'd15890004;
cipher_text[11] = `CIPHERTEXT_WIDTH'd8399794;
cipher_text[12] = `CIPHERTEXT_WIDTH'd1984788;
cipher_text[13] = `CIPHERTEXT_WIDTH'd13751727;
cipher_text[14] = `CIPHERTEXT_WIDTH'd8204486;
cipher_text[15] = `CIPHERTEXT_WIDTH'd7919212;
cipher_text[16] = `CIPHERTEXT_WIDTH'd1297426;
cipher_text[17] = `CIPHERTEXT_WIDTH'd4612046;
cipher_text[18] = `CIPHERTEXT_WIDTH'd16153102;
cipher_text[19] = `CIPHERTEXT_WIDTH'd8484105;
cipher_text[20] = `CIPHERTEXT_WIDTH'd4861269;
cipher_text[21] = `CIPHERTEXT_WIDTH'd10899206;
cipher_text[22] = `CIPHERTEXT_WIDTH'd4965571;
cipher_text[23] = `CIPHERTEXT_WIDTH'd12340285;
cipher_text[24] = `CIPHERTEXT_WIDTH'd7287137;
cipher_text[25] = `CIPHERTEXT_WIDTH'd7513332;
cipher_text[26] = `CIPHERTEXT_WIDTH'd3469086;
cipher_text[27] = `CIPHERTEXT_WIDTH'd4801783;
cipher_text[28] = `CIPHERTEXT_WIDTH'd8149344;
cipher_text[29] = `CIPHERTEXT_WIDTH'd16733343;
cipher_text[30] = `CIPHERTEXT_WIDTH'd1864341;
cipher_text[31] = `CIPHERTEXT_WIDTH'd2032186;
cipher_text[32] = `CIPHERTEXT_WIDTH'd12982499;
cipher_text[33] = `CIPHERTEXT_WIDTH'd7040913;
cipher_text[34] = `CIPHERTEXT_WIDTH'd4639461;
cipher_text[35] = `CIPHERTEXT_WIDTH'd7529733;
cipher_text[36] = `CIPHERTEXT_WIDTH'd9734517;
cipher_text[37] = `CIPHERTEXT_WIDTH'd11738106;
cipher_text[38] = `CIPHERTEXT_WIDTH'd15536660;
cipher_text[39] = `CIPHERTEXT_WIDTH'd971418;
cipher_text[40] = `CIPHERTEXT_WIDTH'd1936329;
cipher_text[41] = `CIPHERTEXT_WIDTH'd9475122;
cipher_text[42] = `CIPHERTEXT_WIDTH'd3220474;
cipher_text[43] = `CIPHERTEXT_WIDTH'd9950409;
cipher_text[44] = `CIPHERTEXT_WIDTH'd3499713;
cipher_text[45] = `CIPHERTEXT_WIDTH'd13544208;
cipher_text[46] = `CIPHERTEXT_WIDTH'd12761332;
cipher_text[47] = `CIPHERTEXT_WIDTH'd6207653;
cipher_text[48] = `CIPHERTEXT_WIDTH'd402004;
cipher_text[49] = `CIPHERTEXT_WIDTH'd14188570;
cipher_text[50] = `CIPHERTEXT_WIDTH'd7972640;
cipher_text[51] = `CIPHERTEXT_WIDTH'd9259777;
cipher_text[52] = `CIPHERTEXT_WIDTH'd7732062;
cipher_text[53] = `CIPHERTEXT_WIDTH'd9772412;
cipher_text[54] = `CIPHERTEXT_WIDTH'd16546570;
cipher_text[55] = `CIPHERTEXT_WIDTH'd5985829;
cipher_text[56] = `CIPHERTEXT_WIDTH'd6935770;
cipher_text[57] = `CIPHERTEXT_WIDTH'd14110667;
cipher_text[58] = `CIPHERTEXT_WIDTH'd13538561;
cipher_text[59] = `CIPHERTEXT_WIDTH'd144899;
cipher_text[60] = `CIPHERTEXT_WIDTH'd5575749;
cipher_text[61] = `CIPHERTEXT_WIDTH'd13594601;
cipher_text[62] = `CIPHERTEXT_WIDTH'd6306020;
cipher_text[63] = `CIPHERTEXT_WIDTH'd6681414;
cipher_text[64] = `CIPHERTEXT_WIDTH'd7506308;
cipher_text[65] = `CIPHERTEXT_WIDTH'd8316373;
cipher_text[66] = `CIPHERTEXT_WIDTH'd2298546;
cipher_text[67] = `CIPHERTEXT_WIDTH'd13304037;
cipher_text[68] = `CIPHERTEXT_WIDTH'd7558333;
cipher_text[69] = `CIPHERTEXT_WIDTH'd3938868;
cipher_text[70] = `CIPHERTEXT_WIDTH'd2648534;
cipher_text[71] = `CIPHERTEXT_WIDTH'd7168632;
cipher_text[72] = `CIPHERTEXT_WIDTH'd5553596;
cipher_text[73] = `CIPHERTEXT_WIDTH'd2963280;
cipher_text[74] = `CIPHERTEXT_WIDTH'd14967156;
cipher_text[75] = `CIPHERTEXT_WIDTH'd15881324;
cipher_text[76] = `CIPHERTEXT_WIDTH'd8371907;
cipher_text[77] = `CIPHERTEXT_WIDTH'd16291234;
cipher_text[78] = `CIPHERTEXT_WIDTH'd7371617;
cipher_text[79] = `CIPHERTEXT_WIDTH'd12870029;
cipher_text[80] = `CIPHERTEXT_WIDTH'd10429900;
cipher_text[81] = `CIPHERTEXT_WIDTH'd11504347;
cipher_text[82] = `CIPHERTEXT_WIDTH'd1641264;
cipher_text[83] = `CIPHERTEXT_WIDTH'd1067081;
cipher_text[84] = `CIPHERTEXT_WIDTH'd2966549;
cipher_text[85] = `CIPHERTEXT_WIDTH'd4997904;
cipher_text[86] = `CIPHERTEXT_WIDTH'd15730220;
cipher_text[87] = `CIPHERTEXT_WIDTH'd3681003;
cipher_text[88] = `CIPHERTEXT_WIDTH'd12870241;
cipher_text[89] = `CIPHERTEXT_WIDTH'd2654099;
cipher_text[90] = `CIPHERTEXT_WIDTH'd9962024;
cipher_text[91] = `CIPHERTEXT_WIDTH'd9269591;
cipher_text[92] = `CIPHERTEXT_WIDTH'd10856943;
cipher_text[93] = `CIPHERTEXT_WIDTH'd15358244;
cipher_text[94] = `CIPHERTEXT_WIDTH'd5852827;
cipher_text[95] = `CIPHERTEXT_WIDTH'd9149768;
cipher_text[96] = `CIPHERTEXT_WIDTH'd7942115;
cipher_text[97] = `CIPHERTEXT_WIDTH'd6579280;
cipher_text[98] = `CIPHERTEXT_WIDTH'd10014749;
cipher_text[99] = `CIPHERTEXT_WIDTH'd4662242;
cipher_text[100] = `CIPHERTEXT_WIDTH'd1952012;
cipher_text[101] = `CIPHERTEXT_WIDTH'd15911655;
cipher_text[102] = `CIPHERTEXT_WIDTH'd4610908;
cipher_text[103] = `CIPHERTEXT_WIDTH'd7345579;
cipher_text[104] = `CIPHERTEXT_WIDTH'd5168715;
cipher_text[105] = `CIPHERTEXT_WIDTH'd12742358;
cipher_text[106] = `CIPHERTEXT_WIDTH'd10095982;
cipher_text[107] = `CIPHERTEXT_WIDTH'd8932750;
cipher_text[108] = `CIPHERTEXT_WIDTH'd1093325;
cipher_text[109] = `CIPHERTEXT_WIDTH'd5627642;
cipher_text[110] = `CIPHERTEXT_WIDTH'd11013560;
cipher_text[111] = `CIPHERTEXT_WIDTH'd10883731;
cipher_text[112] = `CIPHERTEXT_WIDTH'd3256989;
cipher_text[113] = `CIPHERTEXT_WIDTH'd10644372;
cipher_text[114] = `CIPHERTEXT_WIDTH'd5983386;
cipher_text[115] = `CIPHERTEXT_WIDTH'd16503235;
cipher_text[116] = `CIPHERTEXT_WIDTH'd7683638;
cipher_text[117] = `CIPHERTEXT_WIDTH'd7665174;
cipher_text[118] = `CIPHERTEXT_WIDTH'd4898563;
cipher_text[119] = `CIPHERTEXT_WIDTH'd92532;
cipher_text[120] = `CIPHERTEXT_WIDTH'd6216685;
cipher_text[121] = `CIPHERTEXT_WIDTH'd6814350;
cipher_text[122] = `CIPHERTEXT_WIDTH'd1497064;
cipher_text[123] = `CIPHERTEXT_WIDTH'd4354196;
cipher_text[124] = `CIPHERTEXT_WIDTH'd7494186;
cipher_text[125] = `CIPHERTEXT_WIDTH'd15174479;
cipher_text[126] = `CIPHERTEXT_WIDTH'd5343555;
cipher_text[127] = `CIPHERTEXT_WIDTH'd11080676;
cipher_text[128] = `CIPHERTEXT_WIDTH'd884114;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 4;
cipher_text[0] = `CIPHERTEXT_WIDTH'd7439702;
cipher_text[1] = `CIPHERTEXT_WIDTH'd6889072;
cipher_text[2] = `CIPHERTEXT_WIDTH'd11258543;
cipher_text[3] = `CIPHERTEXT_WIDTH'd4392341;
cipher_text[4] = `CIPHERTEXT_WIDTH'd8185952;
cipher_text[5] = `CIPHERTEXT_WIDTH'd7790200;
cipher_text[6] = `CIPHERTEXT_WIDTH'd4391968;
cipher_text[7] = `CIPHERTEXT_WIDTH'd10641757;
cipher_text[8] = `CIPHERTEXT_WIDTH'd6414234;
cipher_text[9] = `CIPHERTEXT_WIDTH'd4351018;
cipher_text[10] = `CIPHERTEXT_WIDTH'd3625121;
cipher_text[11] = `CIPHERTEXT_WIDTH'd2245983;
cipher_text[12] = `CIPHERTEXT_WIDTH'd10268570;
cipher_text[13] = `CIPHERTEXT_WIDTH'd8834627;
cipher_text[14] = `CIPHERTEXT_WIDTH'd279704;
cipher_text[15] = `CIPHERTEXT_WIDTH'd1467895;
cipher_text[16] = `CIPHERTEXT_WIDTH'd3451653;
cipher_text[17] = `CIPHERTEXT_WIDTH'd14936472;
cipher_text[18] = `CIPHERTEXT_WIDTH'd13317804;
cipher_text[19] = `CIPHERTEXT_WIDTH'd7233274;
cipher_text[20] = `CIPHERTEXT_WIDTH'd14076574;
cipher_text[21] = `CIPHERTEXT_WIDTH'd1444122;
cipher_text[22] = `CIPHERTEXT_WIDTH'd10337398;
cipher_text[23] = `CIPHERTEXT_WIDTH'd7576118;
cipher_text[24] = `CIPHERTEXT_WIDTH'd11563972;
cipher_text[25] = `CIPHERTEXT_WIDTH'd5517196;
cipher_text[26] = `CIPHERTEXT_WIDTH'd7926829;
cipher_text[27] = `CIPHERTEXT_WIDTH'd3949142;
cipher_text[28] = `CIPHERTEXT_WIDTH'd12028210;
cipher_text[29] = `CIPHERTEXT_WIDTH'd11883420;
cipher_text[30] = `CIPHERTEXT_WIDTH'd10262812;
cipher_text[31] = `CIPHERTEXT_WIDTH'd1513907;
cipher_text[32] = `CIPHERTEXT_WIDTH'd15764469;
cipher_text[33] = `CIPHERTEXT_WIDTH'd4126783;
cipher_text[34] = `CIPHERTEXT_WIDTH'd5395537;
cipher_text[35] = `CIPHERTEXT_WIDTH'd4526806;
cipher_text[36] = `CIPHERTEXT_WIDTH'd2730477;
cipher_text[37] = `CIPHERTEXT_WIDTH'd1524191;
cipher_text[38] = `CIPHERTEXT_WIDTH'd1585102;
cipher_text[39] = `CIPHERTEXT_WIDTH'd14615966;
cipher_text[40] = `CIPHERTEXT_WIDTH'd7065176;
cipher_text[41] = `CIPHERTEXT_WIDTH'd1316504;
cipher_text[42] = `CIPHERTEXT_WIDTH'd15270042;
cipher_text[43] = `CIPHERTEXT_WIDTH'd15786719;
cipher_text[44] = `CIPHERTEXT_WIDTH'd8836925;
cipher_text[45] = `CIPHERTEXT_WIDTH'd13638117;
cipher_text[46] = `CIPHERTEXT_WIDTH'd12902839;
cipher_text[47] = `CIPHERTEXT_WIDTH'd11207734;
cipher_text[48] = `CIPHERTEXT_WIDTH'd1074559;
cipher_text[49] = `CIPHERTEXT_WIDTH'd2399094;
cipher_text[50] = `CIPHERTEXT_WIDTH'd6586545;
cipher_text[51] = `CIPHERTEXT_WIDTH'd9806412;
cipher_text[52] = `CIPHERTEXT_WIDTH'd3364816;
cipher_text[53] = `CIPHERTEXT_WIDTH'd12140661;
cipher_text[54] = `CIPHERTEXT_WIDTH'd7482630;
cipher_text[55] = `CIPHERTEXT_WIDTH'd8024159;
cipher_text[56] = `CIPHERTEXT_WIDTH'd1362232;
cipher_text[57] = `CIPHERTEXT_WIDTH'd10595586;
cipher_text[58] = `CIPHERTEXT_WIDTH'd9786851;
cipher_text[59] = `CIPHERTEXT_WIDTH'd11749137;
cipher_text[60] = `CIPHERTEXT_WIDTH'd7366569;
cipher_text[61] = `CIPHERTEXT_WIDTH'd1632924;
cipher_text[62] = `CIPHERTEXT_WIDTH'd13356542;
cipher_text[63] = `CIPHERTEXT_WIDTH'd14674251;
cipher_text[64] = `CIPHERTEXT_WIDTH'd4748335;
cipher_text[65] = `CIPHERTEXT_WIDTH'd3156225;
cipher_text[66] = `CIPHERTEXT_WIDTH'd992638;
cipher_text[67] = `CIPHERTEXT_WIDTH'd12193903;
cipher_text[68] = `CIPHERTEXT_WIDTH'd7558553;
cipher_text[69] = `CIPHERTEXT_WIDTH'd14033928;
cipher_text[70] = `CIPHERTEXT_WIDTH'd13422127;
cipher_text[71] = `CIPHERTEXT_WIDTH'd3136916;
cipher_text[72] = `CIPHERTEXT_WIDTH'd15427609;
cipher_text[73] = `CIPHERTEXT_WIDTH'd2006994;
cipher_text[74] = `CIPHERTEXT_WIDTH'd15175386;
cipher_text[75] = `CIPHERTEXT_WIDTH'd1186429;
cipher_text[76] = `CIPHERTEXT_WIDTH'd15968859;
cipher_text[77] = `CIPHERTEXT_WIDTH'd1583766;
cipher_text[78] = `CIPHERTEXT_WIDTH'd7781112;
cipher_text[79] = `CIPHERTEXT_WIDTH'd12509686;
cipher_text[80] = `CIPHERTEXT_WIDTH'd14690497;
cipher_text[81] = `CIPHERTEXT_WIDTH'd4695404;
cipher_text[82] = `CIPHERTEXT_WIDTH'd6504907;
cipher_text[83] = `CIPHERTEXT_WIDTH'd16461633;
cipher_text[84] = `CIPHERTEXT_WIDTH'd2974071;
cipher_text[85] = `CIPHERTEXT_WIDTH'd1030312;
cipher_text[86] = `CIPHERTEXT_WIDTH'd3287029;
cipher_text[87] = `CIPHERTEXT_WIDTH'd6019628;
cipher_text[88] = `CIPHERTEXT_WIDTH'd6707025;
cipher_text[89] = `CIPHERTEXT_WIDTH'd16733795;
cipher_text[90] = `CIPHERTEXT_WIDTH'd12731587;
cipher_text[91] = `CIPHERTEXT_WIDTH'd10056717;
cipher_text[92] = `CIPHERTEXT_WIDTH'd8066319;
cipher_text[93] = `CIPHERTEXT_WIDTH'd4849802;
cipher_text[94] = `CIPHERTEXT_WIDTH'd16510399;
cipher_text[95] = `CIPHERTEXT_WIDTH'd1342084;
cipher_text[96] = `CIPHERTEXT_WIDTH'd16184664;
cipher_text[97] = `CIPHERTEXT_WIDTH'd8576963;
cipher_text[98] = `CIPHERTEXT_WIDTH'd11943488;
cipher_text[99] = `CIPHERTEXT_WIDTH'd6353405;
cipher_text[100] = `CIPHERTEXT_WIDTH'd2114960;
cipher_text[101] = `CIPHERTEXT_WIDTH'd12772101;
cipher_text[102] = `CIPHERTEXT_WIDTH'd2827866;
cipher_text[103] = `CIPHERTEXT_WIDTH'd10437369;
cipher_text[104] = `CIPHERTEXT_WIDTH'd11542576;
cipher_text[105] = `CIPHERTEXT_WIDTH'd8362311;
cipher_text[106] = `CIPHERTEXT_WIDTH'd7525339;
cipher_text[107] = `CIPHERTEXT_WIDTH'd16720467;
cipher_text[108] = `CIPHERTEXT_WIDTH'd3248739;
cipher_text[109] = `CIPHERTEXT_WIDTH'd5367468;
cipher_text[110] = `CIPHERTEXT_WIDTH'd2448198;
cipher_text[111] = `CIPHERTEXT_WIDTH'd5854568;
cipher_text[112] = `CIPHERTEXT_WIDTH'd4740066;
cipher_text[113] = `CIPHERTEXT_WIDTH'd3470005;
cipher_text[114] = `CIPHERTEXT_WIDTH'd11950076;
cipher_text[115] = `CIPHERTEXT_WIDTH'd12041684;
cipher_text[116] = `CIPHERTEXT_WIDTH'd2720006;
cipher_text[117] = `CIPHERTEXT_WIDTH'd2836643;
cipher_text[118] = `CIPHERTEXT_WIDTH'd14362460;
cipher_text[119] = `CIPHERTEXT_WIDTH'd12773169;
cipher_text[120] = `CIPHERTEXT_WIDTH'd14777000;
cipher_text[121] = `CIPHERTEXT_WIDTH'd3666821;
cipher_text[122] = `CIPHERTEXT_WIDTH'd11097230;
cipher_text[123] = `CIPHERTEXT_WIDTH'd4670593;
cipher_text[124] = `CIPHERTEXT_WIDTH'd8514364;
cipher_text[125] = `CIPHERTEXT_WIDTH'd13006372;
cipher_text[126] = `CIPHERTEXT_WIDTH'd2337644;
cipher_text[127] = `CIPHERTEXT_WIDTH'd5537890;
cipher_text[128] = `CIPHERTEXT_WIDTH'd274096;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 5;
cipher_text[0] = `CIPHERTEXT_WIDTH'd15932153;
cipher_text[1] = `CIPHERTEXT_WIDTH'd11420897;
cipher_text[2] = `CIPHERTEXT_WIDTH'd10139537;
cipher_text[3] = `CIPHERTEXT_WIDTH'd1760884;
cipher_text[4] = `CIPHERTEXT_WIDTH'd13316517;
cipher_text[5] = `CIPHERTEXT_WIDTH'd15673978;
cipher_text[6] = `CIPHERTEXT_WIDTH'd10498491;
cipher_text[7] = `CIPHERTEXT_WIDTH'd11183545;
cipher_text[8] = `CIPHERTEXT_WIDTH'd15651585;
cipher_text[9] = `CIPHERTEXT_WIDTH'd2129143;
cipher_text[10] = `CIPHERTEXT_WIDTH'd11196623;
cipher_text[11] = `CIPHERTEXT_WIDTH'd6745021;
cipher_text[12] = `CIPHERTEXT_WIDTH'd14630807;
cipher_text[13] = `CIPHERTEXT_WIDTH'd8300374;
cipher_text[14] = `CIPHERTEXT_WIDTH'd11725080;
cipher_text[15] = `CIPHERTEXT_WIDTH'd7938110;
cipher_text[16] = `CIPHERTEXT_WIDTH'd11879492;
cipher_text[17] = `CIPHERTEXT_WIDTH'd15169031;
cipher_text[18] = `CIPHERTEXT_WIDTH'd14666240;
cipher_text[19] = `CIPHERTEXT_WIDTH'd6582985;
cipher_text[20] = `CIPHERTEXT_WIDTH'd16026225;
cipher_text[21] = `CIPHERTEXT_WIDTH'd14357884;
cipher_text[22] = `CIPHERTEXT_WIDTH'd3711078;
cipher_text[23] = `CIPHERTEXT_WIDTH'd5731168;
cipher_text[24] = `CIPHERTEXT_WIDTH'd11823211;
cipher_text[25] = `CIPHERTEXT_WIDTH'd16380684;
cipher_text[26] = `CIPHERTEXT_WIDTH'd5801162;
cipher_text[27] = `CIPHERTEXT_WIDTH'd2422203;
cipher_text[28] = `CIPHERTEXT_WIDTH'd12496927;
cipher_text[29] = `CIPHERTEXT_WIDTH'd10622610;
cipher_text[30] = `CIPHERTEXT_WIDTH'd12240897;
cipher_text[31] = `CIPHERTEXT_WIDTH'd14561240;
cipher_text[32] = `CIPHERTEXT_WIDTH'd5497086;
cipher_text[33] = `CIPHERTEXT_WIDTH'd16769470;
cipher_text[34] = `CIPHERTEXT_WIDTH'd16041720;
cipher_text[35] = `CIPHERTEXT_WIDTH'd7123548;
cipher_text[36] = `CIPHERTEXT_WIDTH'd6942195;
cipher_text[37] = `CIPHERTEXT_WIDTH'd4143822;
cipher_text[38] = `CIPHERTEXT_WIDTH'd7198550;
cipher_text[39] = `CIPHERTEXT_WIDTH'd4259765;
cipher_text[40] = `CIPHERTEXT_WIDTH'd16045637;
cipher_text[41] = `CIPHERTEXT_WIDTH'd14105986;
cipher_text[42] = `CIPHERTEXT_WIDTH'd6697182;
cipher_text[43] = `CIPHERTEXT_WIDTH'd5169697;
cipher_text[44] = `CIPHERTEXT_WIDTH'd11938855;
cipher_text[45] = `CIPHERTEXT_WIDTH'd7829856;
cipher_text[46] = `CIPHERTEXT_WIDTH'd10521051;
cipher_text[47] = `CIPHERTEXT_WIDTH'd15422057;
cipher_text[48] = `CIPHERTEXT_WIDTH'd10692030;
cipher_text[49] = `CIPHERTEXT_WIDTH'd13494759;
cipher_text[50] = `CIPHERTEXT_WIDTH'd32194;
cipher_text[51] = `CIPHERTEXT_WIDTH'd9688703;
cipher_text[52] = `CIPHERTEXT_WIDTH'd13732925;
cipher_text[53] = `CIPHERTEXT_WIDTH'd13348764;
cipher_text[54] = `CIPHERTEXT_WIDTH'd11567707;
cipher_text[55] = `CIPHERTEXT_WIDTH'd9242514;
cipher_text[56] = `CIPHERTEXT_WIDTH'd7102973;
cipher_text[57] = `CIPHERTEXT_WIDTH'd16675143;
cipher_text[58] = `CIPHERTEXT_WIDTH'd10427861;
cipher_text[59] = `CIPHERTEXT_WIDTH'd6297804;
cipher_text[60] = `CIPHERTEXT_WIDTH'd8674661;
cipher_text[61] = `CIPHERTEXT_WIDTH'd11916320;
cipher_text[62] = `CIPHERTEXT_WIDTH'd13770708;
cipher_text[63] = `CIPHERTEXT_WIDTH'd543427;
cipher_text[64] = `CIPHERTEXT_WIDTH'd10567235;
cipher_text[65] = `CIPHERTEXT_WIDTH'd9973433;
cipher_text[66] = `CIPHERTEXT_WIDTH'd15949657;
cipher_text[67] = `CIPHERTEXT_WIDTH'd7569116;
cipher_text[68] = `CIPHERTEXT_WIDTH'd1503132;
cipher_text[69] = `CIPHERTEXT_WIDTH'd16230299;
cipher_text[70] = `CIPHERTEXT_WIDTH'd6488468;
cipher_text[71] = `CIPHERTEXT_WIDTH'd11981712;
cipher_text[72] = `CIPHERTEXT_WIDTH'd2553636;
cipher_text[73] = `CIPHERTEXT_WIDTH'd2782271;
cipher_text[74] = `CIPHERTEXT_WIDTH'd1407181;
cipher_text[75] = `CIPHERTEXT_WIDTH'd14142224;
cipher_text[76] = `CIPHERTEXT_WIDTH'd8232429;
cipher_text[77] = `CIPHERTEXT_WIDTH'd8727982;
cipher_text[78] = `CIPHERTEXT_WIDTH'd12827636;
cipher_text[79] = `CIPHERTEXT_WIDTH'd10383402;
cipher_text[80] = `CIPHERTEXT_WIDTH'd13632414;
cipher_text[81] = `CIPHERTEXT_WIDTH'd8869943;
cipher_text[82] = `CIPHERTEXT_WIDTH'd15880342;
cipher_text[83] = `CIPHERTEXT_WIDTH'd15215180;
cipher_text[84] = `CIPHERTEXT_WIDTH'd1587390;
cipher_text[85] = `CIPHERTEXT_WIDTH'd11628483;
cipher_text[86] = `CIPHERTEXT_WIDTH'd7879905;
cipher_text[87] = `CIPHERTEXT_WIDTH'd16453897;
cipher_text[88] = `CIPHERTEXT_WIDTH'd2571607;
cipher_text[89] = `CIPHERTEXT_WIDTH'd18320;
cipher_text[90] = `CIPHERTEXT_WIDTH'd12609772;
cipher_text[91] = `CIPHERTEXT_WIDTH'd11011794;
cipher_text[92] = `CIPHERTEXT_WIDTH'd12568963;
cipher_text[93] = `CIPHERTEXT_WIDTH'd5006821;
cipher_text[94] = `CIPHERTEXT_WIDTH'd14494142;
cipher_text[95] = `CIPHERTEXT_WIDTH'd15068740;
cipher_text[96] = `CIPHERTEXT_WIDTH'd11642373;
cipher_text[97] = `CIPHERTEXT_WIDTH'd2510939;
cipher_text[98] = `CIPHERTEXT_WIDTH'd4157501;
cipher_text[99] = `CIPHERTEXT_WIDTH'd12614902;
cipher_text[100] = `CIPHERTEXT_WIDTH'd5697984;
cipher_text[101] = `CIPHERTEXT_WIDTH'd7720744;
cipher_text[102] = `CIPHERTEXT_WIDTH'd11135031;
cipher_text[103] = `CIPHERTEXT_WIDTH'd16055174;
cipher_text[104] = `CIPHERTEXT_WIDTH'd1208471;
cipher_text[105] = `CIPHERTEXT_WIDTH'd6881141;
cipher_text[106] = `CIPHERTEXT_WIDTH'd5414809;
cipher_text[107] = `CIPHERTEXT_WIDTH'd13682138;
cipher_text[108] = `CIPHERTEXT_WIDTH'd13679221;
cipher_text[109] = `CIPHERTEXT_WIDTH'd8945091;
cipher_text[110] = `CIPHERTEXT_WIDTH'd1611008;
cipher_text[111] = `CIPHERTEXT_WIDTH'd11749467;
cipher_text[112] = `CIPHERTEXT_WIDTH'd5945981;
cipher_text[113] = `CIPHERTEXT_WIDTH'd7881115;
cipher_text[114] = `CIPHERTEXT_WIDTH'd6748284;
cipher_text[115] = `CIPHERTEXT_WIDTH'd9890314;
cipher_text[116] = `CIPHERTEXT_WIDTH'd9262105;
cipher_text[117] = `CIPHERTEXT_WIDTH'd10267521;
cipher_text[118] = `CIPHERTEXT_WIDTH'd3708245;
cipher_text[119] = `CIPHERTEXT_WIDTH'd8215239;
cipher_text[120] = `CIPHERTEXT_WIDTH'd4475664;
cipher_text[121] = `CIPHERTEXT_WIDTH'd15034240;
cipher_text[122] = `CIPHERTEXT_WIDTH'd10587198;
cipher_text[123] = `CIPHERTEXT_WIDTH'd8548674;
cipher_text[124] = `CIPHERTEXT_WIDTH'd12355983;
cipher_text[125] = `CIPHERTEXT_WIDTH'd8900036;
cipher_text[126] = `CIPHERTEXT_WIDTH'd12383183;
cipher_text[127] = `CIPHERTEXT_WIDTH'd15388918;
cipher_text[128] = `CIPHERTEXT_WIDTH'd1869366;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 6;
cipher_text[0] = `CIPHERTEXT_WIDTH'd8620265;
cipher_text[1] = `CIPHERTEXT_WIDTH'd6338795;
cipher_text[2] = `CIPHERTEXT_WIDTH'd15624620;
cipher_text[3] = `CIPHERTEXT_WIDTH'd7882506;
cipher_text[4] = `CIPHERTEXT_WIDTH'd12682854;
cipher_text[5] = `CIPHERTEXT_WIDTH'd1034838;
cipher_text[6] = `CIPHERTEXT_WIDTH'd1809027;
cipher_text[7] = `CIPHERTEXT_WIDTH'd6229520;
cipher_text[8] = `CIPHERTEXT_WIDTH'd13331372;
cipher_text[9] = `CIPHERTEXT_WIDTH'd6816255;
cipher_text[10] = `CIPHERTEXT_WIDTH'd9611244;
cipher_text[11] = `CIPHERTEXT_WIDTH'd15799649;
cipher_text[12] = `CIPHERTEXT_WIDTH'd1927943;
cipher_text[13] = `CIPHERTEXT_WIDTH'd13322946;
cipher_text[14] = `CIPHERTEXT_WIDTH'd15860071;
cipher_text[15] = `CIPHERTEXT_WIDTH'd5669111;
cipher_text[16] = `CIPHERTEXT_WIDTH'd2188085;
cipher_text[17] = `CIPHERTEXT_WIDTH'd1265519;
cipher_text[18] = `CIPHERTEXT_WIDTH'd2464147;
cipher_text[19] = `CIPHERTEXT_WIDTH'd3200950;
cipher_text[20] = `CIPHERTEXT_WIDTH'd10583036;
cipher_text[21] = `CIPHERTEXT_WIDTH'd16630578;
cipher_text[22] = `CIPHERTEXT_WIDTH'd16037540;
cipher_text[23] = `CIPHERTEXT_WIDTH'd6853219;
cipher_text[24] = `CIPHERTEXT_WIDTH'd11312344;
cipher_text[25] = `CIPHERTEXT_WIDTH'd6833991;
cipher_text[26] = `CIPHERTEXT_WIDTH'd8914528;
cipher_text[27] = `CIPHERTEXT_WIDTH'd8397104;
cipher_text[28] = `CIPHERTEXT_WIDTH'd13704536;
cipher_text[29] = `CIPHERTEXT_WIDTH'd13514553;
cipher_text[30] = `CIPHERTEXT_WIDTH'd10692286;
cipher_text[31] = `CIPHERTEXT_WIDTH'd39778;
cipher_text[32] = `CIPHERTEXT_WIDTH'd11578983;
cipher_text[33] = `CIPHERTEXT_WIDTH'd11893966;
cipher_text[34] = `CIPHERTEXT_WIDTH'd9792257;
cipher_text[35] = `CIPHERTEXT_WIDTH'd3353830;
cipher_text[36] = `CIPHERTEXT_WIDTH'd1792787;
cipher_text[37] = `CIPHERTEXT_WIDTH'd2898128;
cipher_text[38] = `CIPHERTEXT_WIDTH'd16604911;
cipher_text[39] = `CIPHERTEXT_WIDTH'd756698;
cipher_text[40] = `CIPHERTEXT_WIDTH'd2914205;
cipher_text[41] = `CIPHERTEXT_WIDTH'd2368322;
cipher_text[42] = `CIPHERTEXT_WIDTH'd10268504;
cipher_text[43] = `CIPHERTEXT_WIDTH'd14646591;
cipher_text[44] = `CIPHERTEXT_WIDTH'd2475018;
cipher_text[45] = `CIPHERTEXT_WIDTH'd10896345;
cipher_text[46] = `CIPHERTEXT_WIDTH'd10520610;
cipher_text[47] = `CIPHERTEXT_WIDTH'd9566287;
cipher_text[48] = `CIPHERTEXT_WIDTH'd8260467;
cipher_text[49] = `CIPHERTEXT_WIDTH'd6733030;
cipher_text[50] = `CIPHERTEXT_WIDTH'd13687755;
cipher_text[51] = `CIPHERTEXT_WIDTH'd5755707;
cipher_text[52] = `CIPHERTEXT_WIDTH'd5336228;
cipher_text[53] = `CIPHERTEXT_WIDTH'd3193815;
cipher_text[54] = `CIPHERTEXT_WIDTH'd572643;
cipher_text[55] = `CIPHERTEXT_WIDTH'd11096335;
cipher_text[56] = `CIPHERTEXT_WIDTH'd2501987;
cipher_text[57] = `CIPHERTEXT_WIDTH'd8128867;
cipher_text[58] = `CIPHERTEXT_WIDTH'd16159153;
cipher_text[59] = `CIPHERTEXT_WIDTH'd15279375;
cipher_text[60] = `CIPHERTEXT_WIDTH'd14217600;
cipher_text[61] = `CIPHERTEXT_WIDTH'd16357650;
cipher_text[62] = `CIPHERTEXT_WIDTH'd5212015;
cipher_text[63] = `CIPHERTEXT_WIDTH'd2770108;
cipher_text[64] = `CIPHERTEXT_WIDTH'd10106553;
cipher_text[65] = `CIPHERTEXT_WIDTH'd15916258;
cipher_text[66] = `CIPHERTEXT_WIDTH'd5718210;
cipher_text[67] = `CIPHERTEXT_WIDTH'd15706559;
cipher_text[68] = `CIPHERTEXT_WIDTH'd12215332;
cipher_text[69] = `CIPHERTEXT_WIDTH'd13642780;
cipher_text[70] = `CIPHERTEXT_WIDTH'd9732776;
cipher_text[71] = `CIPHERTEXT_WIDTH'd3605354;
cipher_text[72] = `CIPHERTEXT_WIDTH'd9509573;
cipher_text[73] = `CIPHERTEXT_WIDTH'd7636869;
cipher_text[74] = `CIPHERTEXT_WIDTH'd3430678;
cipher_text[75] = `CIPHERTEXT_WIDTH'd3502760;
cipher_text[76] = `CIPHERTEXT_WIDTH'd14562222;
cipher_text[77] = `CIPHERTEXT_WIDTH'd3196250;
cipher_text[78] = `CIPHERTEXT_WIDTH'd10869314;
cipher_text[79] = `CIPHERTEXT_WIDTH'd14731163;
cipher_text[80] = `CIPHERTEXT_WIDTH'd4930590;
cipher_text[81] = `CIPHERTEXT_WIDTH'd6987518;
cipher_text[82] = `CIPHERTEXT_WIDTH'd10412390;
cipher_text[83] = `CIPHERTEXT_WIDTH'd3468398;
cipher_text[84] = `CIPHERTEXT_WIDTH'd8732347;
cipher_text[85] = `CIPHERTEXT_WIDTH'd569407;
cipher_text[86] = `CIPHERTEXT_WIDTH'd2982548;
cipher_text[87] = `CIPHERTEXT_WIDTH'd14891330;
cipher_text[88] = `CIPHERTEXT_WIDTH'd499793;
cipher_text[89] = `CIPHERTEXT_WIDTH'd3098158;
cipher_text[90] = `CIPHERTEXT_WIDTH'd616661;
cipher_text[91] = `CIPHERTEXT_WIDTH'd16345390;
cipher_text[92] = `CIPHERTEXT_WIDTH'd12796345;
cipher_text[93] = `CIPHERTEXT_WIDTH'd305925;
cipher_text[94] = `CIPHERTEXT_WIDTH'd15727936;
cipher_text[95] = `CIPHERTEXT_WIDTH'd10282951;
cipher_text[96] = `CIPHERTEXT_WIDTH'd16334324;
cipher_text[97] = `CIPHERTEXT_WIDTH'd4205898;
cipher_text[98] = `CIPHERTEXT_WIDTH'd6963182;
cipher_text[99] = `CIPHERTEXT_WIDTH'd1255219;
cipher_text[100] = `CIPHERTEXT_WIDTH'd13924117;
cipher_text[101] = `CIPHERTEXT_WIDTH'd2949246;
cipher_text[102] = `CIPHERTEXT_WIDTH'd6742893;
cipher_text[103] = `CIPHERTEXT_WIDTH'd2753788;
cipher_text[104] = `CIPHERTEXT_WIDTH'd5669172;
cipher_text[105] = `CIPHERTEXT_WIDTH'd5678945;
cipher_text[106] = `CIPHERTEXT_WIDTH'd2349661;
cipher_text[107] = `CIPHERTEXT_WIDTH'd1076401;
cipher_text[108] = `CIPHERTEXT_WIDTH'd11206284;
cipher_text[109] = `CIPHERTEXT_WIDTH'd5160121;
cipher_text[110] = `CIPHERTEXT_WIDTH'd7151934;
cipher_text[111] = `CIPHERTEXT_WIDTH'd10198275;
cipher_text[112] = `CIPHERTEXT_WIDTH'd16168115;
cipher_text[113] = `CIPHERTEXT_WIDTH'd6574024;
cipher_text[114] = `CIPHERTEXT_WIDTH'd243484;
cipher_text[115] = `CIPHERTEXT_WIDTH'd12652099;
cipher_text[116] = `CIPHERTEXT_WIDTH'd5179214;
cipher_text[117] = `CIPHERTEXT_WIDTH'd8519416;
cipher_text[118] = `CIPHERTEXT_WIDTH'd4160329;
cipher_text[119] = `CIPHERTEXT_WIDTH'd3062376;
cipher_text[120] = `CIPHERTEXT_WIDTH'd14696020;
cipher_text[121] = `CIPHERTEXT_WIDTH'd6044578;
cipher_text[122] = `CIPHERTEXT_WIDTH'd14463529;
cipher_text[123] = `CIPHERTEXT_WIDTH'd12887129;
cipher_text[124] = `CIPHERTEXT_WIDTH'd15633156;
cipher_text[125] = `CIPHERTEXT_WIDTH'd13422804;
cipher_text[126] = `CIPHERTEXT_WIDTH'd8036753;
cipher_text[127] = `CIPHERTEXT_WIDTH'd1887962;
cipher_text[128] = `CIPHERTEXT_WIDTH'd12539195;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 7;
cipher_text[0] = `CIPHERTEXT_WIDTH'd7866668;
cipher_text[1] = `CIPHERTEXT_WIDTH'd6780436;
cipher_text[2] = `CIPHERTEXT_WIDTH'd580600;
cipher_text[3] = `CIPHERTEXT_WIDTH'd15653427;
cipher_text[4] = `CIPHERTEXT_WIDTH'd9045358;
cipher_text[5] = `CIPHERTEXT_WIDTH'd14574832;
cipher_text[6] = `CIPHERTEXT_WIDTH'd1947970;
cipher_text[7] = `CIPHERTEXT_WIDTH'd16224876;
cipher_text[8] = `CIPHERTEXT_WIDTH'd15651762;
cipher_text[9] = `CIPHERTEXT_WIDTH'd14709799;
cipher_text[10] = `CIPHERTEXT_WIDTH'd8048567;
cipher_text[11] = `CIPHERTEXT_WIDTH'd5192127;
cipher_text[12] = `CIPHERTEXT_WIDTH'd632223;
cipher_text[13] = `CIPHERTEXT_WIDTH'd10829071;
cipher_text[14] = `CIPHERTEXT_WIDTH'd12320549;
cipher_text[15] = `CIPHERTEXT_WIDTH'd14193512;
cipher_text[16] = `CIPHERTEXT_WIDTH'd7888526;
cipher_text[17] = `CIPHERTEXT_WIDTH'd5548790;
cipher_text[18] = `CIPHERTEXT_WIDTH'd2138966;
cipher_text[19] = `CIPHERTEXT_WIDTH'd3360774;
cipher_text[20] = `CIPHERTEXT_WIDTH'd10542323;
cipher_text[21] = `CIPHERTEXT_WIDTH'd8561984;
cipher_text[22] = `CIPHERTEXT_WIDTH'd4078793;
cipher_text[23] = `CIPHERTEXT_WIDTH'd15892611;
cipher_text[24] = `CIPHERTEXT_WIDTH'd189272;
cipher_text[25] = `CIPHERTEXT_WIDTH'd11290656;
cipher_text[26] = `CIPHERTEXT_WIDTH'd14193988;
cipher_text[27] = `CIPHERTEXT_WIDTH'd10362648;
cipher_text[28] = `CIPHERTEXT_WIDTH'd16042706;
cipher_text[29] = `CIPHERTEXT_WIDTH'd10552529;
cipher_text[30] = `CIPHERTEXT_WIDTH'd16713492;
cipher_text[31] = `CIPHERTEXT_WIDTH'd3502258;
cipher_text[32] = `CIPHERTEXT_WIDTH'd13897251;
cipher_text[33] = `CIPHERTEXT_WIDTH'd11735762;
cipher_text[34] = `CIPHERTEXT_WIDTH'd8756951;
cipher_text[35] = `CIPHERTEXT_WIDTH'd1562456;
cipher_text[36] = `CIPHERTEXT_WIDTH'd2427029;
cipher_text[37] = `CIPHERTEXT_WIDTH'd5744156;
cipher_text[38] = `CIPHERTEXT_WIDTH'd10494023;
cipher_text[39] = `CIPHERTEXT_WIDTH'd5012092;
cipher_text[40] = `CIPHERTEXT_WIDTH'd2054602;
cipher_text[41] = `CIPHERTEXT_WIDTH'd8534028;
cipher_text[42] = `CIPHERTEXT_WIDTH'd1134629;
cipher_text[43] = `CIPHERTEXT_WIDTH'd4957577;
cipher_text[44] = `CIPHERTEXT_WIDTH'd8836443;
cipher_text[45] = `CIPHERTEXT_WIDTH'd7528309;
cipher_text[46] = `CIPHERTEXT_WIDTH'd8425783;
cipher_text[47] = `CIPHERTEXT_WIDTH'd14353027;
cipher_text[48] = `CIPHERTEXT_WIDTH'd8610414;
cipher_text[49] = `CIPHERTEXT_WIDTH'd2570466;
cipher_text[50] = `CIPHERTEXT_WIDTH'd6345004;
cipher_text[51] = `CIPHERTEXT_WIDTH'd10668450;
cipher_text[52] = `CIPHERTEXT_WIDTH'd13956918;
cipher_text[53] = `CIPHERTEXT_WIDTH'd5879547;
cipher_text[54] = `CIPHERTEXT_WIDTH'd846902;
cipher_text[55] = `CIPHERTEXT_WIDTH'd5589849;
cipher_text[56] = `CIPHERTEXT_WIDTH'd5204388;
cipher_text[57] = `CIPHERTEXT_WIDTH'd11324395;
cipher_text[58] = `CIPHERTEXT_WIDTH'd8231475;
cipher_text[59] = `CIPHERTEXT_WIDTH'd903170;
cipher_text[60] = `CIPHERTEXT_WIDTH'd14390250;
cipher_text[61] = `CIPHERTEXT_WIDTH'd114445;
cipher_text[62] = `CIPHERTEXT_WIDTH'd16493927;
cipher_text[63] = `CIPHERTEXT_WIDTH'd260886;
cipher_text[64] = `CIPHERTEXT_WIDTH'd9063052;
cipher_text[65] = `CIPHERTEXT_WIDTH'd6063863;
cipher_text[66] = `CIPHERTEXT_WIDTH'd15868490;
cipher_text[67] = `CIPHERTEXT_WIDTH'd7627019;
cipher_text[68] = `CIPHERTEXT_WIDTH'd6569032;
cipher_text[69] = `CIPHERTEXT_WIDTH'd11093382;
cipher_text[70] = `CIPHERTEXT_WIDTH'd10518254;
cipher_text[71] = `CIPHERTEXT_WIDTH'd13209553;
cipher_text[72] = `CIPHERTEXT_WIDTH'd13074973;
cipher_text[73] = `CIPHERTEXT_WIDTH'd13764690;
cipher_text[74] = `CIPHERTEXT_WIDTH'd8852897;
cipher_text[75] = `CIPHERTEXT_WIDTH'd3088699;
cipher_text[76] = `CIPHERTEXT_WIDTH'd8615796;
cipher_text[77] = `CIPHERTEXT_WIDTH'd4491100;
cipher_text[78] = `CIPHERTEXT_WIDTH'd11799702;
cipher_text[79] = `CIPHERTEXT_WIDTH'd7799858;
cipher_text[80] = `CIPHERTEXT_WIDTH'd13479276;
cipher_text[81] = `CIPHERTEXT_WIDTH'd4424587;
cipher_text[82] = `CIPHERTEXT_WIDTH'd14061613;
cipher_text[83] = `CIPHERTEXT_WIDTH'd6574832;
cipher_text[84] = `CIPHERTEXT_WIDTH'd8355422;
cipher_text[85] = `CIPHERTEXT_WIDTH'd2406671;
cipher_text[86] = `CIPHERTEXT_WIDTH'd9561489;
cipher_text[87] = `CIPHERTEXT_WIDTH'd13104915;
cipher_text[88] = `CIPHERTEXT_WIDTH'd16438936;
cipher_text[89] = `CIPHERTEXT_WIDTH'd3664207;
cipher_text[90] = `CIPHERTEXT_WIDTH'd15129742;
cipher_text[91] = `CIPHERTEXT_WIDTH'd7830282;
cipher_text[92] = `CIPHERTEXT_WIDTH'd14389883;
cipher_text[93] = `CIPHERTEXT_WIDTH'd7299711;
cipher_text[94] = `CIPHERTEXT_WIDTH'd14094949;
cipher_text[95] = `CIPHERTEXT_WIDTH'd13637766;
cipher_text[96] = `CIPHERTEXT_WIDTH'd12915152;
cipher_text[97] = `CIPHERTEXT_WIDTH'd11454242;
cipher_text[98] = `CIPHERTEXT_WIDTH'd2150354;
cipher_text[99] = `CIPHERTEXT_WIDTH'd2133919;
cipher_text[100] = `CIPHERTEXT_WIDTH'd10515195;
cipher_text[101] = `CIPHERTEXT_WIDTH'd861928;
cipher_text[102] = `CIPHERTEXT_WIDTH'd11963858;
cipher_text[103] = `CIPHERTEXT_WIDTH'd14925324;
cipher_text[104] = `CIPHERTEXT_WIDTH'd8324997;
cipher_text[105] = `CIPHERTEXT_WIDTH'd1888504;
cipher_text[106] = `CIPHERTEXT_WIDTH'd16413035;
cipher_text[107] = `CIPHERTEXT_WIDTH'd939831;
cipher_text[108] = `CIPHERTEXT_WIDTH'd1184832;
cipher_text[109] = `CIPHERTEXT_WIDTH'd10542886;
cipher_text[110] = `CIPHERTEXT_WIDTH'd9854393;
cipher_text[111] = `CIPHERTEXT_WIDTH'd13566930;
cipher_text[112] = `CIPHERTEXT_WIDTH'd721290;
cipher_text[113] = `CIPHERTEXT_WIDTH'd6535431;
cipher_text[114] = `CIPHERTEXT_WIDTH'd3624187;
cipher_text[115] = `CIPHERTEXT_WIDTH'd8876737;
cipher_text[116] = `CIPHERTEXT_WIDTH'd16508346;
cipher_text[117] = `CIPHERTEXT_WIDTH'd6591653;
cipher_text[118] = `CIPHERTEXT_WIDTH'd13419485;
cipher_text[119] = `CIPHERTEXT_WIDTH'd15964699;
cipher_text[120] = `CIPHERTEXT_WIDTH'd9335639;
cipher_text[121] = `CIPHERTEXT_WIDTH'd1703220;
cipher_text[122] = `CIPHERTEXT_WIDTH'd3087797;
cipher_text[123] = `CIPHERTEXT_WIDTH'd6137122;
cipher_text[124] = `CIPHERTEXT_WIDTH'd2907241;
cipher_text[125] = `CIPHERTEXT_WIDTH'd12775837;
cipher_text[126] = `CIPHERTEXT_WIDTH'd2831088;
cipher_text[127] = `CIPHERTEXT_WIDTH'd10431220;
cipher_text[128] = `CIPHERTEXT_WIDTH'd13845428;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 8;
cipher_text[0] = `CIPHERTEXT_WIDTH'd2855433;
cipher_text[1] = `CIPHERTEXT_WIDTH'd2386746;
cipher_text[2] = `CIPHERTEXT_WIDTH'd10174669;
cipher_text[3] = `CIPHERTEXT_WIDTH'd12162553;
cipher_text[4] = `CIPHERTEXT_WIDTH'd8072006;
cipher_text[5] = `CIPHERTEXT_WIDTH'd1281140;
cipher_text[6] = `CIPHERTEXT_WIDTH'd717973;
cipher_text[7] = `CIPHERTEXT_WIDTH'd9152774;
cipher_text[8] = `CIPHERTEXT_WIDTH'd11658808;
cipher_text[9] = `CIPHERTEXT_WIDTH'd11736930;
cipher_text[10] = `CIPHERTEXT_WIDTH'd5470220;
cipher_text[11] = `CIPHERTEXT_WIDTH'd6822558;
cipher_text[12] = `CIPHERTEXT_WIDTH'd11718025;
cipher_text[13] = `CIPHERTEXT_WIDTH'd7320634;
cipher_text[14] = `CIPHERTEXT_WIDTH'd5116170;
cipher_text[15] = `CIPHERTEXT_WIDTH'd16229770;
cipher_text[16] = `CIPHERTEXT_WIDTH'd4144101;
cipher_text[17] = `CIPHERTEXT_WIDTH'd10244046;
cipher_text[18] = `CIPHERTEXT_WIDTH'd4705846;
cipher_text[19] = `CIPHERTEXT_WIDTH'd3249977;
cipher_text[20] = `CIPHERTEXT_WIDTH'd15938063;
cipher_text[21] = `CIPHERTEXT_WIDTH'd13306791;
cipher_text[22] = `CIPHERTEXT_WIDTH'd8836285;
cipher_text[23] = `CIPHERTEXT_WIDTH'd10701603;
cipher_text[24] = `CIPHERTEXT_WIDTH'd8014754;
cipher_text[25] = `CIPHERTEXT_WIDTH'd3557585;
cipher_text[26] = `CIPHERTEXT_WIDTH'd14158833;
cipher_text[27] = `CIPHERTEXT_WIDTH'd13214096;
cipher_text[28] = `CIPHERTEXT_WIDTH'd9335531;
cipher_text[29] = `CIPHERTEXT_WIDTH'd12358404;
cipher_text[30] = `CIPHERTEXT_WIDTH'd8260321;
cipher_text[31] = `CIPHERTEXT_WIDTH'd14508786;
cipher_text[32] = `CIPHERTEXT_WIDTH'd2433532;
cipher_text[33] = `CIPHERTEXT_WIDTH'd11129368;
cipher_text[34] = `CIPHERTEXT_WIDTH'd16603722;
cipher_text[35] = `CIPHERTEXT_WIDTH'd7508324;
cipher_text[36] = `CIPHERTEXT_WIDTH'd2162850;
cipher_text[37] = `CIPHERTEXT_WIDTH'd1452033;
cipher_text[38] = `CIPHERTEXT_WIDTH'd10153718;
cipher_text[39] = `CIPHERTEXT_WIDTH'd9368533;
cipher_text[40] = `CIPHERTEXT_WIDTH'd196091;
cipher_text[41] = `CIPHERTEXT_WIDTH'd13338509;
cipher_text[42] = `CIPHERTEXT_WIDTH'd14736418;
cipher_text[43] = `CIPHERTEXT_WIDTH'd7363437;
cipher_text[44] = `CIPHERTEXT_WIDTH'd16218129;
cipher_text[45] = `CIPHERTEXT_WIDTH'd10960396;
cipher_text[46] = `CIPHERTEXT_WIDTH'd12290002;
cipher_text[47] = `CIPHERTEXT_WIDTH'd3171872;
cipher_text[48] = `CIPHERTEXT_WIDTH'd11854663;
cipher_text[49] = `CIPHERTEXT_WIDTH'd12357066;
cipher_text[50] = `CIPHERTEXT_WIDTH'd11697893;
cipher_text[51] = `CIPHERTEXT_WIDTH'd2616853;
cipher_text[52] = `CIPHERTEXT_WIDTH'd5064103;
cipher_text[53] = `CIPHERTEXT_WIDTH'd13514230;
cipher_text[54] = `CIPHERTEXT_WIDTH'd8907181;
cipher_text[55] = `CIPHERTEXT_WIDTH'd2673645;
cipher_text[56] = `CIPHERTEXT_WIDTH'd15302690;
cipher_text[57] = `CIPHERTEXT_WIDTH'd5737550;
cipher_text[58] = `CIPHERTEXT_WIDTH'd2099174;
cipher_text[59] = `CIPHERTEXT_WIDTH'd1520357;
cipher_text[60] = `CIPHERTEXT_WIDTH'd6706024;
cipher_text[61] = `CIPHERTEXT_WIDTH'd1311654;
cipher_text[62] = `CIPHERTEXT_WIDTH'd610307;
cipher_text[63] = `CIPHERTEXT_WIDTH'd9130676;
cipher_text[64] = `CIPHERTEXT_WIDTH'd15267990;
cipher_text[65] = `CIPHERTEXT_WIDTH'd9979443;
cipher_text[66] = `CIPHERTEXT_WIDTH'd15345607;
cipher_text[67] = `CIPHERTEXT_WIDTH'd397994;
cipher_text[68] = `CIPHERTEXT_WIDTH'd14784652;
cipher_text[69] = `CIPHERTEXT_WIDTH'd5160117;
cipher_text[70] = `CIPHERTEXT_WIDTH'd11478707;
cipher_text[71] = `CIPHERTEXT_WIDTH'd8817270;
cipher_text[72] = `CIPHERTEXT_WIDTH'd7188385;
cipher_text[73] = `CIPHERTEXT_WIDTH'd14340107;
cipher_text[74] = `CIPHERTEXT_WIDTH'd16061900;
cipher_text[75] = `CIPHERTEXT_WIDTH'd2168503;
cipher_text[76] = `CIPHERTEXT_WIDTH'd4613953;
cipher_text[77] = `CIPHERTEXT_WIDTH'd2292350;
cipher_text[78] = `CIPHERTEXT_WIDTH'd2115721;
cipher_text[79] = `CIPHERTEXT_WIDTH'd10384432;
cipher_text[80] = `CIPHERTEXT_WIDTH'd7137729;
cipher_text[81] = `CIPHERTEXT_WIDTH'd15285480;
cipher_text[82] = `CIPHERTEXT_WIDTH'd11333410;
cipher_text[83] = `CIPHERTEXT_WIDTH'd14980184;
cipher_text[84] = `CIPHERTEXT_WIDTH'd3795105;
cipher_text[85] = `CIPHERTEXT_WIDTH'd9090617;
cipher_text[86] = `CIPHERTEXT_WIDTH'd2037605;
cipher_text[87] = `CIPHERTEXT_WIDTH'd6739773;
cipher_text[88] = `CIPHERTEXT_WIDTH'd8547970;
cipher_text[89] = `CIPHERTEXT_WIDTH'd15285408;
cipher_text[90] = `CIPHERTEXT_WIDTH'd7772617;
cipher_text[91] = `CIPHERTEXT_WIDTH'd9180664;
cipher_text[92] = `CIPHERTEXT_WIDTH'd10028358;
cipher_text[93] = `CIPHERTEXT_WIDTH'd5463608;
cipher_text[94] = `CIPHERTEXT_WIDTH'd15090846;
cipher_text[95] = `CIPHERTEXT_WIDTH'd5261655;
cipher_text[96] = `CIPHERTEXT_WIDTH'd5395539;
cipher_text[97] = `CIPHERTEXT_WIDTH'd7715785;
cipher_text[98] = `CIPHERTEXT_WIDTH'd3858614;
cipher_text[99] = `CIPHERTEXT_WIDTH'd8358890;
cipher_text[100] = `CIPHERTEXT_WIDTH'd14245016;
cipher_text[101] = `CIPHERTEXT_WIDTH'd3630032;
cipher_text[102] = `CIPHERTEXT_WIDTH'd10789253;
cipher_text[103] = `CIPHERTEXT_WIDTH'd10414696;
cipher_text[104] = `CIPHERTEXT_WIDTH'd8667764;
cipher_text[105] = `CIPHERTEXT_WIDTH'd14315320;
cipher_text[106] = `CIPHERTEXT_WIDTH'd9838591;
cipher_text[107] = `CIPHERTEXT_WIDTH'd7087985;
cipher_text[108] = `CIPHERTEXT_WIDTH'd5735098;
cipher_text[109] = `CIPHERTEXT_WIDTH'd10357685;
cipher_text[110] = `CIPHERTEXT_WIDTH'd1708224;
cipher_text[111] = `CIPHERTEXT_WIDTH'd13746286;
cipher_text[112] = `CIPHERTEXT_WIDTH'd4849361;
cipher_text[113] = `CIPHERTEXT_WIDTH'd12433775;
cipher_text[114] = `CIPHERTEXT_WIDTH'd1698272;
cipher_text[115] = `CIPHERTEXT_WIDTH'd3361625;
cipher_text[116] = `CIPHERTEXT_WIDTH'd6911437;
cipher_text[117] = `CIPHERTEXT_WIDTH'd16172512;
cipher_text[118] = `CIPHERTEXT_WIDTH'd436944;
cipher_text[119] = `CIPHERTEXT_WIDTH'd11163339;
cipher_text[120] = `CIPHERTEXT_WIDTH'd13850485;
cipher_text[121] = `CIPHERTEXT_WIDTH'd12480615;
cipher_text[122] = `CIPHERTEXT_WIDTH'd24211;
cipher_text[123] = `CIPHERTEXT_WIDTH'd11491830;
cipher_text[124] = `CIPHERTEXT_WIDTH'd6404832;
cipher_text[125] = `CIPHERTEXT_WIDTH'd6502579;
cipher_text[126] = `CIPHERTEXT_WIDTH'd16265500;
cipher_text[127] = `CIPHERTEXT_WIDTH'd14976988;
cipher_text[128] = `CIPHERTEXT_WIDTH'd10762781;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 9;
cipher_text[0] = `CIPHERTEXT_WIDTH'd3000560;
cipher_text[1] = `CIPHERTEXT_WIDTH'd12584540;
cipher_text[2] = `CIPHERTEXT_WIDTH'd851662;
cipher_text[3] = `CIPHERTEXT_WIDTH'd267525;
cipher_text[4] = `CIPHERTEXT_WIDTH'd13904809;
cipher_text[5] = `CIPHERTEXT_WIDTH'd8409841;
cipher_text[6] = `CIPHERTEXT_WIDTH'd6784986;
cipher_text[7] = `CIPHERTEXT_WIDTH'd1258106;
cipher_text[8] = `CIPHERTEXT_WIDTH'd15992154;
cipher_text[9] = `CIPHERTEXT_WIDTH'd5756711;
cipher_text[10] = `CIPHERTEXT_WIDTH'd16748981;
cipher_text[11] = `CIPHERTEXT_WIDTH'd30492;
cipher_text[12] = `CIPHERTEXT_WIDTH'd8902542;
cipher_text[13] = `CIPHERTEXT_WIDTH'd10172117;
cipher_text[14] = `CIPHERTEXT_WIDTH'd9081957;
cipher_text[15] = `CIPHERTEXT_WIDTH'd3065560;
cipher_text[16] = `CIPHERTEXT_WIDTH'd9679899;
cipher_text[17] = `CIPHERTEXT_WIDTH'd6549552;
cipher_text[18] = `CIPHERTEXT_WIDTH'd15702641;
cipher_text[19] = `CIPHERTEXT_WIDTH'd10474230;
cipher_text[20] = `CIPHERTEXT_WIDTH'd7222702;
cipher_text[21] = `CIPHERTEXT_WIDTH'd366530;
cipher_text[22] = `CIPHERTEXT_WIDTH'd5954546;
cipher_text[23] = `CIPHERTEXT_WIDTH'd3533069;
cipher_text[24] = `CIPHERTEXT_WIDTH'd7240951;
cipher_text[25] = `CIPHERTEXT_WIDTH'd7073404;
cipher_text[26] = `CIPHERTEXT_WIDTH'd8449148;
cipher_text[27] = `CIPHERTEXT_WIDTH'd8238595;
cipher_text[28] = `CIPHERTEXT_WIDTH'd8089136;
cipher_text[29] = `CIPHERTEXT_WIDTH'd13097066;
cipher_text[30] = `CIPHERTEXT_WIDTH'd4348430;
cipher_text[31] = `CIPHERTEXT_WIDTH'd11136878;
cipher_text[32] = `CIPHERTEXT_WIDTH'd10801697;
cipher_text[33] = `CIPHERTEXT_WIDTH'd15190730;
cipher_text[34] = `CIPHERTEXT_WIDTH'd3055597;
cipher_text[35] = `CIPHERTEXT_WIDTH'd9627206;
cipher_text[36] = `CIPHERTEXT_WIDTH'd4255115;
cipher_text[37] = `CIPHERTEXT_WIDTH'd6051170;
cipher_text[38] = `CIPHERTEXT_WIDTH'd8486173;
cipher_text[39] = `CIPHERTEXT_WIDTH'd13106574;
cipher_text[40] = `CIPHERTEXT_WIDTH'd11417958;
cipher_text[41] = `CIPHERTEXT_WIDTH'd9869993;
cipher_text[42] = `CIPHERTEXT_WIDTH'd11143919;
cipher_text[43] = `CIPHERTEXT_WIDTH'd14704792;
cipher_text[44] = `CIPHERTEXT_WIDTH'd224291;
cipher_text[45] = `CIPHERTEXT_WIDTH'd4599844;
cipher_text[46] = `CIPHERTEXT_WIDTH'd13321604;
cipher_text[47] = `CIPHERTEXT_WIDTH'd15511717;
cipher_text[48] = `CIPHERTEXT_WIDTH'd6632920;
cipher_text[49] = `CIPHERTEXT_WIDTH'd14177274;
cipher_text[50] = `CIPHERTEXT_WIDTH'd8831336;
cipher_text[51] = `CIPHERTEXT_WIDTH'd4896207;
cipher_text[52] = `CIPHERTEXT_WIDTH'd10793984;
cipher_text[53] = `CIPHERTEXT_WIDTH'd13691933;
cipher_text[54] = `CIPHERTEXT_WIDTH'd9028110;
cipher_text[55] = `CIPHERTEXT_WIDTH'd7855116;
cipher_text[56] = `CIPHERTEXT_WIDTH'd5392056;
cipher_text[57] = `CIPHERTEXT_WIDTH'd12929726;
cipher_text[58] = `CIPHERTEXT_WIDTH'd6453868;
cipher_text[59] = `CIPHERTEXT_WIDTH'd14838949;
cipher_text[60] = `CIPHERTEXT_WIDTH'd8677065;
cipher_text[61] = `CIPHERTEXT_WIDTH'd5959282;
cipher_text[62] = `CIPHERTEXT_WIDTH'd4352442;
cipher_text[63] = `CIPHERTEXT_WIDTH'd7397773;
cipher_text[64] = `CIPHERTEXT_WIDTH'd864046;
cipher_text[65] = `CIPHERTEXT_WIDTH'd10086646;
cipher_text[66] = `CIPHERTEXT_WIDTH'd101746;
cipher_text[67] = `CIPHERTEXT_WIDTH'd7694887;
cipher_text[68] = `CIPHERTEXT_WIDTH'd9075110;
cipher_text[69] = `CIPHERTEXT_WIDTH'd14288602;
cipher_text[70] = `CIPHERTEXT_WIDTH'd8993370;
cipher_text[71] = `CIPHERTEXT_WIDTH'd368867;
cipher_text[72] = `CIPHERTEXT_WIDTH'd6299159;
cipher_text[73] = `CIPHERTEXT_WIDTH'd13686916;
cipher_text[74] = `CIPHERTEXT_WIDTH'd16160144;
cipher_text[75] = `CIPHERTEXT_WIDTH'd8980995;
cipher_text[76] = `CIPHERTEXT_WIDTH'd3008309;
cipher_text[77] = `CIPHERTEXT_WIDTH'd16164548;
cipher_text[78] = `CIPHERTEXT_WIDTH'd15936240;
cipher_text[79] = `CIPHERTEXT_WIDTH'd16678709;
cipher_text[80] = `CIPHERTEXT_WIDTH'd12896578;
cipher_text[81] = `CIPHERTEXT_WIDTH'd2180704;
cipher_text[82] = `CIPHERTEXT_WIDTH'd548506;
cipher_text[83] = `CIPHERTEXT_WIDTH'd9510064;
cipher_text[84] = `CIPHERTEXT_WIDTH'd1672252;
cipher_text[85] = `CIPHERTEXT_WIDTH'd12393297;
cipher_text[86] = `CIPHERTEXT_WIDTH'd3752869;
cipher_text[87] = `CIPHERTEXT_WIDTH'd6329379;
cipher_text[88] = `CIPHERTEXT_WIDTH'd705430;
cipher_text[89] = `CIPHERTEXT_WIDTH'd13124244;
cipher_text[90] = `CIPHERTEXT_WIDTH'd4011458;
cipher_text[91] = `CIPHERTEXT_WIDTH'd3704581;
cipher_text[92] = `CIPHERTEXT_WIDTH'd8796316;
cipher_text[93] = `CIPHERTEXT_WIDTH'd15319015;
cipher_text[94] = `CIPHERTEXT_WIDTH'd217310;
cipher_text[95] = `CIPHERTEXT_WIDTH'd7304702;
cipher_text[96] = `CIPHERTEXT_WIDTH'd4862272;
cipher_text[97] = `CIPHERTEXT_WIDTH'd3617996;
cipher_text[98] = `CIPHERTEXT_WIDTH'd3160744;
cipher_text[99] = `CIPHERTEXT_WIDTH'd1805040;
cipher_text[100] = `CIPHERTEXT_WIDTH'd6206729;
cipher_text[101] = `CIPHERTEXT_WIDTH'd15207860;
cipher_text[102] = `CIPHERTEXT_WIDTH'd8692455;
cipher_text[103] = `CIPHERTEXT_WIDTH'd10331544;
cipher_text[104] = `CIPHERTEXT_WIDTH'd9681872;
cipher_text[105] = `CIPHERTEXT_WIDTH'd7914765;
cipher_text[106] = `CIPHERTEXT_WIDTH'd13594782;
cipher_text[107] = `CIPHERTEXT_WIDTH'd488702;
cipher_text[108] = `CIPHERTEXT_WIDTH'd10982711;
cipher_text[109] = `CIPHERTEXT_WIDTH'd8486525;
cipher_text[110] = `CIPHERTEXT_WIDTH'd6051499;
cipher_text[111] = `CIPHERTEXT_WIDTH'd10101633;
cipher_text[112] = `CIPHERTEXT_WIDTH'd7161808;
cipher_text[113] = `CIPHERTEXT_WIDTH'd10007484;
cipher_text[114] = `CIPHERTEXT_WIDTH'd6856274;
cipher_text[115] = `CIPHERTEXT_WIDTH'd2148843;
cipher_text[116] = `CIPHERTEXT_WIDTH'd7645700;
cipher_text[117] = `CIPHERTEXT_WIDTH'd2766529;
cipher_text[118] = `CIPHERTEXT_WIDTH'd10296673;
cipher_text[119] = `CIPHERTEXT_WIDTH'd7223411;
cipher_text[120] = `CIPHERTEXT_WIDTH'd466428;
cipher_text[121] = `CIPHERTEXT_WIDTH'd10694002;
cipher_text[122] = `CIPHERTEXT_WIDTH'd9463247;
cipher_text[123] = `CIPHERTEXT_WIDTH'd1997546;
cipher_text[124] = `CIPHERTEXT_WIDTH'd14736709;
cipher_text[125] = `CIPHERTEXT_WIDTH'd15567540;
cipher_text[126] = `CIPHERTEXT_WIDTH'd2143867;
cipher_text[127] = `CIPHERTEXT_WIDTH'd3771938;
cipher_text[128] = `CIPHERTEXT_WIDTH'd3710942;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 10;
cipher_text[0] = `CIPHERTEXT_WIDTH'd2928967;
cipher_text[1] = `CIPHERTEXT_WIDTH'd14053596;
cipher_text[2] = `CIPHERTEXT_WIDTH'd12863323;
cipher_text[3] = `CIPHERTEXT_WIDTH'd3207872;
cipher_text[4] = `CIPHERTEXT_WIDTH'd8806408;
cipher_text[5] = `CIPHERTEXT_WIDTH'd9101215;
cipher_text[6] = `CIPHERTEXT_WIDTH'd14233152;
cipher_text[7] = `CIPHERTEXT_WIDTH'd5808654;
cipher_text[8] = `CIPHERTEXT_WIDTH'd15702052;
cipher_text[9] = `CIPHERTEXT_WIDTH'd13062982;
cipher_text[10] = `CIPHERTEXT_WIDTH'd5626291;
cipher_text[11] = `CIPHERTEXT_WIDTH'd773121;
cipher_text[12] = `CIPHERTEXT_WIDTH'd3223119;
cipher_text[13] = `CIPHERTEXT_WIDTH'd1738371;
cipher_text[14] = `CIPHERTEXT_WIDTH'd6459574;
cipher_text[15] = `CIPHERTEXT_WIDTH'd7095483;
cipher_text[16] = `CIPHERTEXT_WIDTH'd666336;
cipher_text[17] = `CIPHERTEXT_WIDTH'd5695087;
cipher_text[18] = `CIPHERTEXT_WIDTH'd10716836;
cipher_text[19] = `CIPHERTEXT_WIDTH'd2340013;
cipher_text[20] = `CIPHERTEXT_WIDTH'd13568811;
cipher_text[21] = `CIPHERTEXT_WIDTH'd6719354;
cipher_text[22] = `CIPHERTEXT_WIDTH'd15607412;
cipher_text[23] = `CIPHERTEXT_WIDTH'd10773167;
cipher_text[24] = `CIPHERTEXT_WIDTH'd3985174;
cipher_text[25] = `CIPHERTEXT_WIDTH'd3575870;
cipher_text[26] = `CIPHERTEXT_WIDTH'd12593549;
cipher_text[27] = `CIPHERTEXT_WIDTH'd10753985;
cipher_text[28] = `CIPHERTEXT_WIDTH'd8375332;
cipher_text[29] = `CIPHERTEXT_WIDTH'd10603755;
cipher_text[30] = `CIPHERTEXT_WIDTH'd8035899;
cipher_text[31] = `CIPHERTEXT_WIDTH'd8181759;
cipher_text[32] = `CIPHERTEXT_WIDTH'd11977237;
cipher_text[33] = `CIPHERTEXT_WIDTH'd13724081;
cipher_text[34] = `CIPHERTEXT_WIDTH'd10916623;
cipher_text[35] = `CIPHERTEXT_WIDTH'd15339110;
cipher_text[36] = `CIPHERTEXT_WIDTH'd3409243;
cipher_text[37] = `CIPHERTEXT_WIDTH'd13866097;
cipher_text[38] = `CIPHERTEXT_WIDTH'd3866449;
cipher_text[39] = `CIPHERTEXT_WIDTH'd471676;
cipher_text[40] = `CIPHERTEXT_WIDTH'd3201292;
cipher_text[41] = `CIPHERTEXT_WIDTH'd9055952;
cipher_text[42] = `CIPHERTEXT_WIDTH'd7136798;
cipher_text[43] = `CIPHERTEXT_WIDTH'd14763141;
cipher_text[44] = `CIPHERTEXT_WIDTH'd5667612;
cipher_text[45] = `CIPHERTEXT_WIDTH'd370534;
cipher_text[46] = `CIPHERTEXT_WIDTH'd9557555;
cipher_text[47] = `CIPHERTEXT_WIDTH'd9069541;
cipher_text[48] = `CIPHERTEXT_WIDTH'd2756511;
cipher_text[49] = `CIPHERTEXT_WIDTH'd11212647;
cipher_text[50] = `CIPHERTEXT_WIDTH'd9361579;
cipher_text[51] = `CIPHERTEXT_WIDTH'd9707131;
cipher_text[52] = `CIPHERTEXT_WIDTH'd976179;
cipher_text[53] = `CIPHERTEXT_WIDTH'd2914556;
cipher_text[54] = `CIPHERTEXT_WIDTH'd5024778;
cipher_text[55] = `CIPHERTEXT_WIDTH'd3441024;
cipher_text[56] = `CIPHERTEXT_WIDTH'd11966175;
cipher_text[57] = `CIPHERTEXT_WIDTH'd16237920;
cipher_text[58] = `CIPHERTEXT_WIDTH'd8976670;
cipher_text[59] = `CIPHERTEXT_WIDTH'd10240037;
cipher_text[60] = `CIPHERTEXT_WIDTH'd7433581;
cipher_text[61] = `CIPHERTEXT_WIDTH'd10845280;
cipher_text[62] = `CIPHERTEXT_WIDTH'd29413;
cipher_text[63] = `CIPHERTEXT_WIDTH'd14964736;
cipher_text[64] = `CIPHERTEXT_WIDTH'd7783445;
cipher_text[65] = `CIPHERTEXT_WIDTH'd12081758;
cipher_text[66] = `CIPHERTEXT_WIDTH'd12636694;
cipher_text[67] = `CIPHERTEXT_WIDTH'd12935283;
cipher_text[68] = `CIPHERTEXT_WIDTH'd11340569;
cipher_text[69] = `CIPHERTEXT_WIDTH'd3465760;
cipher_text[70] = `CIPHERTEXT_WIDTH'd7676490;
cipher_text[71] = `CIPHERTEXT_WIDTH'd5040525;
cipher_text[72] = `CIPHERTEXT_WIDTH'd3533784;
cipher_text[73] = `CIPHERTEXT_WIDTH'd1719093;
cipher_text[74] = `CIPHERTEXT_WIDTH'd13628503;
cipher_text[75] = `CIPHERTEXT_WIDTH'd12830234;
cipher_text[76] = `CIPHERTEXT_WIDTH'd2843743;
cipher_text[77] = `CIPHERTEXT_WIDTH'd8395336;
cipher_text[78] = `CIPHERTEXT_WIDTH'd6391441;
cipher_text[79] = `CIPHERTEXT_WIDTH'd4782549;
cipher_text[80] = `CIPHERTEXT_WIDTH'd12400841;
cipher_text[81] = `CIPHERTEXT_WIDTH'd11145435;
cipher_text[82] = `CIPHERTEXT_WIDTH'd2986140;
cipher_text[83] = `CIPHERTEXT_WIDTH'd13806142;
cipher_text[84] = `CIPHERTEXT_WIDTH'd11180774;
cipher_text[85] = `CIPHERTEXT_WIDTH'd8664363;
cipher_text[86] = `CIPHERTEXT_WIDTH'd6254050;
cipher_text[87] = `CIPHERTEXT_WIDTH'd7377335;
cipher_text[88] = `CIPHERTEXT_WIDTH'd1334899;
cipher_text[89] = `CIPHERTEXT_WIDTH'd16072290;
cipher_text[90] = `CIPHERTEXT_WIDTH'd12366233;
cipher_text[91] = `CIPHERTEXT_WIDTH'd11884742;
cipher_text[92] = `CIPHERTEXT_WIDTH'd1114530;
cipher_text[93] = `CIPHERTEXT_WIDTH'd2212265;
cipher_text[94] = `CIPHERTEXT_WIDTH'd3383109;
cipher_text[95] = `CIPHERTEXT_WIDTH'd10127759;
cipher_text[96] = `CIPHERTEXT_WIDTH'd11662025;
cipher_text[97] = `CIPHERTEXT_WIDTH'd12207322;
cipher_text[98] = `CIPHERTEXT_WIDTH'd6354710;
cipher_text[99] = `CIPHERTEXT_WIDTH'd12571705;
cipher_text[100] = `CIPHERTEXT_WIDTH'd5719459;
cipher_text[101] = `CIPHERTEXT_WIDTH'd14666383;
cipher_text[102] = `CIPHERTEXT_WIDTH'd16528381;
cipher_text[103] = `CIPHERTEXT_WIDTH'd15716549;
cipher_text[104] = `CIPHERTEXT_WIDTH'd8484159;
cipher_text[105] = `CIPHERTEXT_WIDTH'd13374710;
cipher_text[106] = `CIPHERTEXT_WIDTH'd205915;
cipher_text[107] = `CIPHERTEXT_WIDTH'd10261482;
cipher_text[108] = `CIPHERTEXT_WIDTH'd12350132;
cipher_text[109] = `CIPHERTEXT_WIDTH'd2093289;
cipher_text[110] = `CIPHERTEXT_WIDTH'd6646085;
cipher_text[111] = `CIPHERTEXT_WIDTH'd5375687;
cipher_text[112] = `CIPHERTEXT_WIDTH'd3598830;
cipher_text[113] = `CIPHERTEXT_WIDTH'd6342701;
cipher_text[114] = `CIPHERTEXT_WIDTH'd13716005;
cipher_text[115] = `CIPHERTEXT_WIDTH'd8858610;
cipher_text[116] = `CIPHERTEXT_WIDTH'd8269410;
cipher_text[117] = `CIPHERTEXT_WIDTH'd5679881;
cipher_text[118] = `CIPHERTEXT_WIDTH'd747033;
cipher_text[119] = `CIPHERTEXT_WIDTH'd4074193;
cipher_text[120] = `CIPHERTEXT_WIDTH'd2505338;
cipher_text[121] = `CIPHERTEXT_WIDTH'd10536153;
cipher_text[122] = `CIPHERTEXT_WIDTH'd4259194;
cipher_text[123] = `CIPHERTEXT_WIDTH'd6192302;
cipher_text[124] = `CIPHERTEXT_WIDTH'd7894183;
cipher_text[125] = `CIPHERTEXT_WIDTH'd8812853;
cipher_text[126] = `CIPHERTEXT_WIDTH'd9695330;
cipher_text[127] = `CIPHERTEXT_WIDTH'd1024636;
cipher_text[128] = `CIPHERTEXT_WIDTH'd16452423;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 11;
cipher_text[0] = `CIPHERTEXT_WIDTH'd5166185;
cipher_text[1] = `CIPHERTEXT_WIDTH'd14550792;
cipher_text[2] = `CIPHERTEXT_WIDTH'd10534278;
cipher_text[3] = `CIPHERTEXT_WIDTH'd23751;
cipher_text[4] = `CIPHERTEXT_WIDTH'd11506085;
cipher_text[5] = `CIPHERTEXT_WIDTH'd15556178;
cipher_text[6] = `CIPHERTEXT_WIDTH'd11288866;
cipher_text[7] = `CIPHERTEXT_WIDTH'd14383244;
cipher_text[8] = `CIPHERTEXT_WIDTH'd16441272;
cipher_text[9] = `CIPHERTEXT_WIDTH'd7128957;
cipher_text[10] = `CIPHERTEXT_WIDTH'd13755455;
cipher_text[11] = `CIPHERTEXT_WIDTH'd4013887;
cipher_text[12] = `CIPHERTEXT_WIDTH'd1580898;
cipher_text[13] = `CIPHERTEXT_WIDTH'd2905291;
cipher_text[14] = `CIPHERTEXT_WIDTH'd13318339;
cipher_text[15] = `CIPHERTEXT_WIDTH'd8083399;
cipher_text[16] = `CIPHERTEXT_WIDTH'd1137817;
cipher_text[17] = `CIPHERTEXT_WIDTH'd13787170;
cipher_text[18] = `CIPHERTEXT_WIDTH'd269258;
cipher_text[19] = `CIPHERTEXT_WIDTH'd7079764;
cipher_text[20] = `CIPHERTEXT_WIDTH'd13668424;
cipher_text[21] = `CIPHERTEXT_WIDTH'd1581035;
cipher_text[22] = `CIPHERTEXT_WIDTH'd10142756;
cipher_text[23] = `CIPHERTEXT_WIDTH'd4401328;
cipher_text[24] = `CIPHERTEXT_WIDTH'd7486617;
cipher_text[25] = `CIPHERTEXT_WIDTH'd808587;
cipher_text[26] = `CIPHERTEXT_WIDTH'd941177;
cipher_text[27] = `CIPHERTEXT_WIDTH'd2264930;
cipher_text[28] = `CIPHERTEXT_WIDTH'd3167465;
cipher_text[29] = `CIPHERTEXT_WIDTH'd8937494;
cipher_text[30] = `CIPHERTEXT_WIDTH'd14681000;
cipher_text[31] = `CIPHERTEXT_WIDTH'd3848017;
cipher_text[32] = `CIPHERTEXT_WIDTH'd12168288;
cipher_text[33] = `CIPHERTEXT_WIDTH'd16562272;
cipher_text[34] = `CIPHERTEXT_WIDTH'd13673975;
cipher_text[35] = `CIPHERTEXT_WIDTH'd12422922;
cipher_text[36] = `CIPHERTEXT_WIDTH'd6752645;
cipher_text[37] = `CIPHERTEXT_WIDTH'd10325937;
cipher_text[38] = `CIPHERTEXT_WIDTH'd10731201;
cipher_text[39] = `CIPHERTEXT_WIDTH'd3900425;
cipher_text[40] = `CIPHERTEXT_WIDTH'd8681141;
cipher_text[41] = `CIPHERTEXT_WIDTH'd550047;
cipher_text[42] = `CIPHERTEXT_WIDTH'd8663378;
cipher_text[43] = `CIPHERTEXT_WIDTH'd873376;
cipher_text[44] = `CIPHERTEXT_WIDTH'd14522835;
cipher_text[45] = `CIPHERTEXT_WIDTH'd2014042;
cipher_text[46] = `CIPHERTEXT_WIDTH'd946026;
cipher_text[47] = `CIPHERTEXT_WIDTH'd5654861;
cipher_text[48] = `CIPHERTEXT_WIDTH'd15668299;
cipher_text[49] = `CIPHERTEXT_WIDTH'd13451436;
cipher_text[50] = `CIPHERTEXT_WIDTH'd3844772;
cipher_text[51] = `CIPHERTEXT_WIDTH'd14456258;
cipher_text[52] = `CIPHERTEXT_WIDTH'd15710056;
cipher_text[53] = `CIPHERTEXT_WIDTH'd6572331;
cipher_text[54] = `CIPHERTEXT_WIDTH'd15929779;
cipher_text[55] = `CIPHERTEXT_WIDTH'd3199463;
cipher_text[56] = `CIPHERTEXT_WIDTH'd12935121;
cipher_text[57] = `CIPHERTEXT_WIDTH'd12618805;
cipher_text[58] = `CIPHERTEXT_WIDTH'd15962754;
cipher_text[59] = `CIPHERTEXT_WIDTH'd13030734;
cipher_text[60] = `CIPHERTEXT_WIDTH'd14970927;
cipher_text[61] = `CIPHERTEXT_WIDTH'd12793277;
cipher_text[62] = `CIPHERTEXT_WIDTH'd6077505;
cipher_text[63] = `CIPHERTEXT_WIDTH'd12635197;
cipher_text[64] = `CIPHERTEXT_WIDTH'd283292;
cipher_text[65] = `CIPHERTEXT_WIDTH'd3203109;
cipher_text[66] = `CIPHERTEXT_WIDTH'd5798633;
cipher_text[67] = `CIPHERTEXT_WIDTH'd10033839;
cipher_text[68] = `CIPHERTEXT_WIDTH'd8117353;
cipher_text[69] = `CIPHERTEXT_WIDTH'd4421074;
cipher_text[70] = `CIPHERTEXT_WIDTH'd13427046;
cipher_text[71] = `CIPHERTEXT_WIDTH'd14800611;
cipher_text[72] = `CIPHERTEXT_WIDTH'd5700297;
cipher_text[73] = `CIPHERTEXT_WIDTH'd9484738;
cipher_text[74] = `CIPHERTEXT_WIDTH'd9418514;
cipher_text[75] = `CIPHERTEXT_WIDTH'd13308077;
cipher_text[76] = `CIPHERTEXT_WIDTH'd5424090;
cipher_text[77] = `CIPHERTEXT_WIDTH'd12450415;
cipher_text[78] = `CIPHERTEXT_WIDTH'd12401555;
cipher_text[79] = `CIPHERTEXT_WIDTH'd1562704;
cipher_text[80] = `CIPHERTEXT_WIDTH'd6849553;
cipher_text[81] = `CIPHERTEXT_WIDTH'd10283711;
cipher_text[82] = `CIPHERTEXT_WIDTH'd10228038;
cipher_text[83] = `CIPHERTEXT_WIDTH'd15848502;
cipher_text[84] = `CIPHERTEXT_WIDTH'd4941313;
cipher_text[85] = `CIPHERTEXT_WIDTH'd1907263;
cipher_text[86] = `CIPHERTEXT_WIDTH'd9144574;
cipher_text[87] = `CIPHERTEXT_WIDTH'd8585414;
cipher_text[88] = `CIPHERTEXT_WIDTH'd8147604;
cipher_text[89] = `CIPHERTEXT_WIDTH'd5229276;
cipher_text[90] = `CIPHERTEXT_WIDTH'd8120411;
cipher_text[91] = `CIPHERTEXT_WIDTH'd3660135;
cipher_text[92] = `CIPHERTEXT_WIDTH'd13539333;
cipher_text[93] = `CIPHERTEXT_WIDTH'd2985654;
cipher_text[94] = `CIPHERTEXT_WIDTH'd2216825;
cipher_text[95] = `CIPHERTEXT_WIDTH'd13542071;
cipher_text[96] = `CIPHERTEXT_WIDTH'd12870545;
cipher_text[97] = `CIPHERTEXT_WIDTH'd7898384;
cipher_text[98] = `CIPHERTEXT_WIDTH'd9942599;
cipher_text[99] = `CIPHERTEXT_WIDTH'd3524818;
cipher_text[100] = `CIPHERTEXT_WIDTH'd8502716;
cipher_text[101] = `CIPHERTEXT_WIDTH'd8918002;
cipher_text[102] = `CIPHERTEXT_WIDTH'd6219358;
cipher_text[103] = `CIPHERTEXT_WIDTH'd4656006;
cipher_text[104] = `CIPHERTEXT_WIDTH'd4883471;
cipher_text[105] = `CIPHERTEXT_WIDTH'd5638308;
cipher_text[106] = `CIPHERTEXT_WIDTH'd3449930;
cipher_text[107] = `CIPHERTEXT_WIDTH'd97129;
cipher_text[108] = `CIPHERTEXT_WIDTH'd2073406;
cipher_text[109] = `CIPHERTEXT_WIDTH'd16744758;
cipher_text[110] = `CIPHERTEXT_WIDTH'd7755603;
cipher_text[111] = `CIPHERTEXT_WIDTH'd6997134;
cipher_text[112] = `CIPHERTEXT_WIDTH'd4539736;
cipher_text[113] = `CIPHERTEXT_WIDTH'd11903040;
cipher_text[114] = `CIPHERTEXT_WIDTH'd1577258;
cipher_text[115] = `CIPHERTEXT_WIDTH'd15636423;
cipher_text[116] = `CIPHERTEXT_WIDTH'd16644238;
cipher_text[117] = `CIPHERTEXT_WIDTH'd9786276;
cipher_text[118] = `CIPHERTEXT_WIDTH'd579104;
cipher_text[119] = `CIPHERTEXT_WIDTH'd974798;
cipher_text[120] = `CIPHERTEXT_WIDTH'd14396508;
cipher_text[121] = `CIPHERTEXT_WIDTH'd620538;
cipher_text[122] = `CIPHERTEXT_WIDTH'd2181061;
cipher_text[123] = `CIPHERTEXT_WIDTH'd4498807;
cipher_text[124] = `CIPHERTEXT_WIDTH'd4675820;
cipher_text[125] = `CIPHERTEXT_WIDTH'd12973840;
cipher_text[126] = `CIPHERTEXT_WIDTH'd15932434;
cipher_text[127] = `CIPHERTEXT_WIDTH'd5253834;
cipher_text[128] = `CIPHERTEXT_WIDTH'd2617828;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 12;
cipher_text[0] = `CIPHERTEXT_WIDTH'd4029023;
cipher_text[1] = `CIPHERTEXT_WIDTH'd4174754;
cipher_text[2] = `CIPHERTEXT_WIDTH'd7229182;
cipher_text[3] = `CIPHERTEXT_WIDTH'd6442056;
cipher_text[4] = `CIPHERTEXT_WIDTH'd12669115;
cipher_text[5] = `CIPHERTEXT_WIDTH'd1251337;
cipher_text[6] = `CIPHERTEXT_WIDTH'd474771;
cipher_text[7] = `CIPHERTEXT_WIDTH'd14762555;
cipher_text[8] = `CIPHERTEXT_WIDTH'd9830034;
cipher_text[9] = `CIPHERTEXT_WIDTH'd13410996;
cipher_text[10] = `CIPHERTEXT_WIDTH'd15511045;
cipher_text[11] = `CIPHERTEXT_WIDTH'd6579089;
cipher_text[12] = `CIPHERTEXT_WIDTH'd5761106;
cipher_text[13] = `CIPHERTEXT_WIDTH'd9129496;
cipher_text[14] = `CIPHERTEXT_WIDTH'd3788857;
cipher_text[15] = `CIPHERTEXT_WIDTH'd6325798;
cipher_text[16] = `CIPHERTEXT_WIDTH'd9597153;
cipher_text[17] = `CIPHERTEXT_WIDTH'd3393251;
cipher_text[18] = `CIPHERTEXT_WIDTH'd7893191;
cipher_text[19] = `CIPHERTEXT_WIDTH'd3314582;
cipher_text[20] = `CIPHERTEXT_WIDTH'd4736972;
cipher_text[21] = `CIPHERTEXT_WIDTH'd10840524;
cipher_text[22] = `CIPHERTEXT_WIDTH'd5748996;
cipher_text[23] = `CIPHERTEXT_WIDTH'd13558820;
cipher_text[24] = `CIPHERTEXT_WIDTH'd9919954;
cipher_text[25] = `CIPHERTEXT_WIDTH'd10389916;
cipher_text[26] = `CIPHERTEXT_WIDTH'd6500124;
cipher_text[27] = `CIPHERTEXT_WIDTH'd3791638;
cipher_text[28] = `CIPHERTEXT_WIDTH'd15824543;
cipher_text[29] = `CIPHERTEXT_WIDTH'd9145263;
cipher_text[30] = `CIPHERTEXT_WIDTH'd4739701;
cipher_text[31] = `CIPHERTEXT_WIDTH'd2821667;
cipher_text[32] = `CIPHERTEXT_WIDTH'd6441329;
cipher_text[33] = `CIPHERTEXT_WIDTH'd3528559;
cipher_text[34] = `CIPHERTEXT_WIDTH'd9019502;
cipher_text[35] = `CIPHERTEXT_WIDTH'd5078090;
cipher_text[36] = `CIPHERTEXT_WIDTH'd12488037;
cipher_text[37] = `CIPHERTEXT_WIDTH'd15909450;
cipher_text[38] = `CIPHERTEXT_WIDTH'd13557458;
cipher_text[39] = `CIPHERTEXT_WIDTH'd373239;
cipher_text[40] = `CIPHERTEXT_WIDTH'd11681792;
cipher_text[41] = `CIPHERTEXT_WIDTH'd4940486;
cipher_text[42] = `CIPHERTEXT_WIDTH'd16126756;
cipher_text[43] = `CIPHERTEXT_WIDTH'd11770679;
cipher_text[44] = `CIPHERTEXT_WIDTH'd3957034;
cipher_text[45] = `CIPHERTEXT_WIDTH'd8951533;
cipher_text[46] = `CIPHERTEXT_WIDTH'd4508432;
cipher_text[47] = `CIPHERTEXT_WIDTH'd8275908;
cipher_text[48] = `CIPHERTEXT_WIDTH'd12801074;
cipher_text[49] = `CIPHERTEXT_WIDTH'd3585263;
cipher_text[50] = `CIPHERTEXT_WIDTH'd9830344;
cipher_text[51] = `CIPHERTEXT_WIDTH'd5513851;
cipher_text[52] = `CIPHERTEXT_WIDTH'd2539088;
cipher_text[53] = `CIPHERTEXT_WIDTH'd2243035;
cipher_text[54] = `CIPHERTEXT_WIDTH'd14909514;
cipher_text[55] = `CIPHERTEXT_WIDTH'd1346761;
cipher_text[56] = `CIPHERTEXT_WIDTH'd2721839;
cipher_text[57] = `CIPHERTEXT_WIDTH'd12125211;
cipher_text[58] = `CIPHERTEXT_WIDTH'd1935800;
cipher_text[59] = `CIPHERTEXT_WIDTH'd2643411;
cipher_text[60] = `CIPHERTEXT_WIDTH'd16728253;
cipher_text[61] = `CIPHERTEXT_WIDTH'd13124370;
cipher_text[62] = `CIPHERTEXT_WIDTH'd1452350;
cipher_text[63] = `CIPHERTEXT_WIDTH'd11663189;
cipher_text[64] = `CIPHERTEXT_WIDTH'd10202864;
cipher_text[65] = `CIPHERTEXT_WIDTH'd10667356;
cipher_text[66] = `CIPHERTEXT_WIDTH'd7409606;
cipher_text[67] = `CIPHERTEXT_WIDTH'd16578522;
cipher_text[68] = `CIPHERTEXT_WIDTH'd16328102;
cipher_text[69] = `CIPHERTEXT_WIDTH'd13791824;
cipher_text[70] = `CIPHERTEXT_WIDTH'd2477901;
cipher_text[71] = `CIPHERTEXT_WIDTH'd3201912;
cipher_text[72] = `CIPHERTEXT_WIDTH'd9736036;
cipher_text[73] = `CIPHERTEXT_WIDTH'd1352273;
cipher_text[74] = `CIPHERTEXT_WIDTH'd15446028;
cipher_text[75] = `CIPHERTEXT_WIDTH'd8128282;
cipher_text[76] = `CIPHERTEXT_WIDTH'd6165734;
cipher_text[77] = `CIPHERTEXT_WIDTH'd15204773;
cipher_text[78] = `CIPHERTEXT_WIDTH'd12598445;
cipher_text[79] = `CIPHERTEXT_WIDTH'd8699590;
cipher_text[80] = `CIPHERTEXT_WIDTH'd8170613;
cipher_text[81] = `CIPHERTEXT_WIDTH'd8350265;
cipher_text[82] = `CIPHERTEXT_WIDTH'd12784950;
cipher_text[83] = `CIPHERTEXT_WIDTH'd6349870;
cipher_text[84] = `CIPHERTEXT_WIDTH'd6267356;
cipher_text[85] = `CIPHERTEXT_WIDTH'd12920579;
cipher_text[86] = `CIPHERTEXT_WIDTH'd15582941;
cipher_text[87] = `CIPHERTEXT_WIDTH'd14943667;
cipher_text[88] = `CIPHERTEXT_WIDTH'd6931993;
cipher_text[89] = `CIPHERTEXT_WIDTH'd10350537;
cipher_text[90] = `CIPHERTEXT_WIDTH'd10462597;
cipher_text[91] = `CIPHERTEXT_WIDTH'd13376378;
cipher_text[92] = `CIPHERTEXT_WIDTH'd4057376;
cipher_text[93] = `CIPHERTEXT_WIDTH'd15411144;
cipher_text[94] = `CIPHERTEXT_WIDTH'd1882135;
cipher_text[95] = `CIPHERTEXT_WIDTH'd2739953;
cipher_text[96] = `CIPHERTEXT_WIDTH'd6436925;
cipher_text[97] = `CIPHERTEXT_WIDTH'd13448291;
cipher_text[98] = `CIPHERTEXT_WIDTH'd2943931;
cipher_text[99] = `CIPHERTEXT_WIDTH'd4429089;
cipher_text[100] = `CIPHERTEXT_WIDTH'd14892011;
cipher_text[101] = `CIPHERTEXT_WIDTH'd11162958;
cipher_text[102] = `CIPHERTEXT_WIDTH'd6573952;
cipher_text[103] = `CIPHERTEXT_WIDTH'd9736859;
cipher_text[104] = `CIPHERTEXT_WIDTH'd1053418;
cipher_text[105] = `CIPHERTEXT_WIDTH'd2404061;
cipher_text[106] = `CIPHERTEXT_WIDTH'd11704506;
cipher_text[107] = `CIPHERTEXT_WIDTH'd3993893;
cipher_text[108] = `CIPHERTEXT_WIDTH'd4626620;
cipher_text[109] = `CIPHERTEXT_WIDTH'd15894543;
cipher_text[110] = `CIPHERTEXT_WIDTH'd1247481;
cipher_text[111] = `CIPHERTEXT_WIDTH'd12618524;
cipher_text[112] = `CIPHERTEXT_WIDTH'd8745106;
cipher_text[113] = `CIPHERTEXT_WIDTH'd14737309;
cipher_text[114] = `CIPHERTEXT_WIDTH'd1158841;
cipher_text[115] = `CIPHERTEXT_WIDTH'd9535951;
cipher_text[116] = `CIPHERTEXT_WIDTH'd4149196;
cipher_text[117] = `CIPHERTEXT_WIDTH'd9869365;
cipher_text[118] = `CIPHERTEXT_WIDTH'd10183136;
cipher_text[119] = `CIPHERTEXT_WIDTH'd12492158;
cipher_text[120] = `CIPHERTEXT_WIDTH'd9335230;
cipher_text[121] = `CIPHERTEXT_WIDTH'd12945812;
cipher_text[122] = `CIPHERTEXT_WIDTH'd8522267;
cipher_text[123] = `CIPHERTEXT_WIDTH'd1247490;
cipher_text[124] = `CIPHERTEXT_WIDTH'd12080155;
cipher_text[125] = `CIPHERTEXT_WIDTH'd9250743;
cipher_text[126] = `CIPHERTEXT_WIDTH'd4322486;
cipher_text[127] = `CIPHERTEXT_WIDTH'd9054670;
cipher_text[128] = `CIPHERTEXT_WIDTH'd2364444;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 13;
cipher_text[0] = `CIPHERTEXT_WIDTH'd4299312;
cipher_text[1] = `CIPHERTEXT_WIDTH'd2873440;
cipher_text[2] = `CIPHERTEXT_WIDTH'd580673;
cipher_text[3] = `CIPHERTEXT_WIDTH'd3157039;
cipher_text[4] = `CIPHERTEXT_WIDTH'd3698995;
cipher_text[5] = `CIPHERTEXT_WIDTH'd4389225;
cipher_text[6] = `CIPHERTEXT_WIDTH'd4642555;
cipher_text[7] = `CIPHERTEXT_WIDTH'd6736436;
cipher_text[8] = `CIPHERTEXT_WIDTH'd10385374;
cipher_text[9] = `CIPHERTEXT_WIDTH'd11571782;
cipher_text[10] = `CIPHERTEXT_WIDTH'd4352331;
cipher_text[11] = `CIPHERTEXT_WIDTH'd15792687;
cipher_text[12] = `CIPHERTEXT_WIDTH'd5943495;
cipher_text[13] = `CIPHERTEXT_WIDTH'd4910934;
cipher_text[14] = `CIPHERTEXT_WIDTH'd9410215;
cipher_text[15] = `CIPHERTEXT_WIDTH'd1710534;
cipher_text[16] = `CIPHERTEXT_WIDTH'd10375151;
cipher_text[17] = `CIPHERTEXT_WIDTH'd13642285;
cipher_text[18] = `CIPHERTEXT_WIDTH'd9853142;
cipher_text[19] = `CIPHERTEXT_WIDTH'd14081762;
cipher_text[20] = `CIPHERTEXT_WIDTH'd10177776;
cipher_text[21] = `CIPHERTEXT_WIDTH'd15800488;
cipher_text[22] = `CIPHERTEXT_WIDTH'd6372164;
cipher_text[23] = `CIPHERTEXT_WIDTH'd1858731;
cipher_text[24] = `CIPHERTEXT_WIDTH'd3988495;
cipher_text[25] = `CIPHERTEXT_WIDTH'd1690651;
cipher_text[26] = `CIPHERTEXT_WIDTH'd6364399;
cipher_text[27] = `CIPHERTEXT_WIDTH'd2675275;
cipher_text[28] = `CIPHERTEXT_WIDTH'd10009739;
cipher_text[29] = `CIPHERTEXT_WIDTH'd1108952;
cipher_text[30] = `CIPHERTEXT_WIDTH'd2463579;
cipher_text[31] = `CIPHERTEXT_WIDTH'd9886260;
cipher_text[32] = `CIPHERTEXT_WIDTH'd3567832;
cipher_text[33] = `CIPHERTEXT_WIDTH'd14290176;
cipher_text[34] = `CIPHERTEXT_WIDTH'd15707312;
cipher_text[35] = `CIPHERTEXT_WIDTH'd14844214;
cipher_text[36] = `CIPHERTEXT_WIDTH'd4821296;
cipher_text[37] = `CIPHERTEXT_WIDTH'd1863771;
cipher_text[38] = `CIPHERTEXT_WIDTH'd10930777;
cipher_text[39] = `CIPHERTEXT_WIDTH'd3054865;
cipher_text[40] = `CIPHERTEXT_WIDTH'd8492878;
cipher_text[41] = `CIPHERTEXT_WIDTH'd623064;
cipher_text[42] = `CIPHERTEXT_WIDTH'd4359905;
cipher_text[43] = `CIPHERTEXT_WIDTH'd1586723;
cipher_text[44] = `CIPHERTEXT_WIDTH'd5954456;
cipher_text[45] = `CIPHERTEXT_WIDTH'd16433316;
cipher_text[46] = `CIPHERTEXT_WIDTH'd11175574;
cipher_text[47] = `CIPHERTEXT_WIDTH'd7374931;
cipher_text[48] = `CIPHERTEXT_WIDTH'd16677476;
cipher_text[49] = `CIPHERTEXT_WIDTH'd10526185;
cipher_text[50] = `CIPHERTEXT_WIDTH'd5311763;
cipher_text[51] = `CIPHERTEXT_WIDTH'd1800922;
cipher_text[52] = `CIPHERTEXT_WIDTH'd8123476;
cipher_text[53] = `CIPHERTEXT_WIDTH'd14671392;
cipher_text[54] = `CIPHERTEXT_WIDTH'd16147906;
cipher_text[55] = `CIPHERTEXT_WIDTH'd11277429;
cipher_text[56] = `CIPHERTEXT_WIDTH'd9361216;
cipher_text[57] = `CIPHERTEXT_WIDTH'd14205439;
cipher_text[58] = `CIPHERTEXT_WIDTH'd15983500;
cipher_text[59] = `CIPHERTEXT_WIDTH'd14311993;
cipher_text[60] = `CIPHERTEXT_WIDTH'd3246797;
cipher_text[61] = `CIPHERTEXT_WIDTH'd12958839;
cipher_text[62] = `CIPHERTEXT_WIDTH'd3651125;
cipher_text[63] = `CIPHERTEXT_WIDTH'd8703292;
cipher_text[64] = `CIPHERTEXT_WIDTH'd14495190;
cipher_text[65] = `CIPHERTEXT_WIDTH'd2479892;
cipher_text[66] = `CIPHERTEXT_WIDTH'd7327851;
cipher_text[67] = `CIPHERTEXT_WIDTH'd2643063;
cipher_text[68] = `CIPHERTEXT_WIDTH'd10461671;
cipher_text[69] = `CIPHERTEXT_WIDTH'd12618784;
cipher_text[70] = `CIPHERTEXT_WIDTH'd10184633;
cipher_text[71] = `CIPHERTEXT_WIDTH'd14997952;
cipher_text[72] = `CIPHERTEXT_WIDTH'd11293775;
cipher_text[73] = `CIPHERTEXT_WIDTH'd4159420;
cipher_text[74] = `CIPHERTEXT_WIDTH'd13871915;
cipher_text[75] = `CIPHERTEXT_WIDTH'd4890008;
cipher_text[76] = `CIPHERTEXT_WIDTH'd8662547;
cipher_text[77] = `CIPHERTEXT_WIDTH'd14625230;
cipher_text[78] = `CIPHERTEXT_WIDTH'd4689432;
cipher_text[79] = `CIPHERTEXT_WIDTH'd12171941;
cipher_text[80] = `CIPHERTEXT_WIDTH'd7150988;
cipher_text[81] = `CIPHERTEXT_WIDTH'd5679961;
cipher_text[82] = `CIPHERTEXT_WIDTH'd10087239;
cipher_text[83] = `CIPHERTEXT_WIDTH'd13056278;
cipher_text[84] = `CIPHERTEXT_WIDTH'd9712028;
cipher_text[85] = `CIPHERTEXT_WIDTH'd5688004;
cipher_text[86] = `CIPHERTEXT_WIDTH'd11628157;
cipher_text[87] = `CIPHERTEXT_WIDTH'd5194515;
cipher_text[88] = `CIPHERTEXT_WIDTH'd11563618;
cipher_text[89] = `CIPHERTEXT_WIDTH'd15544817;
cipher_text[90] = `CIPHERTEXT_WIDTH'd7338839;
cipher_text[91] = `CIPHERTEXT_WIDTH'd16247194;
cipher_text[92] = `CIPHERTEXT_WIDTH'd15472295;
cipher_text[93] = `CIPHERTEXT_WIDTH'd10389103;
cipher_text[94] = `CIPHERTEXT_WIDTH'd5102630;
cipher_text[95] = `CIPHERTEXT_WIDTH'd4363867;
cipher_text[96] = `CIPHERTEXT_WIDTH'd13556058;
cipher_text[97] = `CIPHERTEXT_WIDTH'd13687005;
cipher_text[98] = `CIPHERTEXT_WIDTH'd1614712;
cipher_text[99] = `CIPHERTEXT_WIDTH'd6565353;
cipher_text[100] = `CIPHERTEXT_WIDTH'd2038249;
cipher_text[101] = `CIPHERTEXT_WIDTH'd4669945;
cipher_text[102] = `CIPHERTEXT_WIDTH'd7932329;
cipher_text[103] = `CIPHERTEXT_WIDTH'd10650312;
cipher_text[104] = `CIPHERTEXT_WIDTH'd2311332;
cipher_text[105] = `CIPHERTEXT_WIDTH'd2044940;
cipher_text[106] = `CIPHERTEXT_WIDTH'd13388270;
cipher_text[107] = `CIPHERTEXT_WIDTH'd8179003;
cipher_text[108] = `CIPHERTEXT_WIDTH'd9622906;
cipher_text[109] = `CIPHERTEXT_WIDTH'd406074;
cipher_text[110] = `CIPHERTEXT_WIDTH'd10270466;
cipher_text[111] = `CIPHERTEXT_WIDTH'd5440247;
cipher_text[112] = `CIPHERTEXT_WIDTH'd12652423;
cipher_text[113] = `CIPHERTEXT_WIDTH'd2128014;
cipher_text[114] = `CIPHERTEXT_WIDTH'd3073054;
cipher_text[115] = `CIPHERTEXT_WIDTH'd4080232;
cipher_text[116] = `CIPHERTEXT_WIDTH'd10552689;
cipher_text[117] = `CIPHERTEXT_WIDTH'd16680322;
cipher_text[118] = `CIPHERTEXT_WIDTH'd5954024;
cipher_text[119] = `CIPHERTEXT_WIDTH'd9685757;
cipher_text[120] = `CIPHERTEXT_WIDTH'd5331063;
cipher_text[121] = `CIPHERTEXT_WIDTH'd9551345;
cipher_text[122] = `CIPHERTEXT_WIDTH'd11687822;
cipher_text[123] = `CIPHERTEXT_WIDTH'd2367212;
cipher_text[124] = `CIPHERTEXT_WIDTH'd9626250;
cipher_text[125] = `CIPHERTEXT_WIDTH'd9400719;
cipher_text[126] = `CIPHERTEXT_WIDTH'd12567088;
cipher_text[127] = `CIPHERTEXT_WIDTH'd3329317;
cipher_text[128] = `CIPHERTEXT_WIDTH'd6189549;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 14;
cipher_text[0] = `CIPHERTEXT_WIDTH'd5422332;
cipher_text[1] = `CIPHERTEXT_WIDTH'd16268011;
cipher_text[2] = `CIPHERTEXT_WIDTH'd8527441;
cipher_text[3] = `CIPHERTEXT_WIDTH'd16207404;
cipher_text[4] = `CIPHERTEXT_WIDTH'd15447252;
cipher_text[5] = `CIPHERTEXT_WIDTH'd12765058;
cipher_text[6] = `CIPHERTEXT_WIDTH'd14166256;
cipher_text[7] = `CIPHERTEXT_WIDTH'd9407060;
cipher_text[8] = `CIPHERTEXT_WIDTH'd15351158;
cipher_text[9] = `CIPHERTEXT_WIDTH'd14447249;
cipher_text[10] = `CIPHERTEXT_WIDTH'd10585313;
cipher_text[11] = `CIPHERTEXT_WIDTH'd8460545;
cipher_text[12] = `CIPHERTEXT_WIDTH'd16159316;
cipher_text[13] = `CIPHERTEXT_WIDTH'd16397086;
cipher_text[14] = `CIPHERTEXT_WIDTH'd1257026;
cipher_text[15] = `CIPHERTEXT_WIDTH'd12322187;
cipher_text[16] = `CIPHERTEXT_WIDTH'd12487672;
cipher_text[17] = `CIPHERTEXT_WIDTH'd12766344;
cipher_text[18] = `CIPHERTEXT_WIDTH'd7790986;
cipher_text[19] = `CIPHERTEXT_WIDTH'd16238155;
cipher_text[20] = `CIPHERTEXT_WIDTH'd15168655;
cipher_text[21] = `CIPHERTEXT_WIDTH'd8619043;
cipher_text[22] = `CIPHERTEXT_WIDTH'd3852706;
cipher_text[23] = `CIPHERTEXT_WIDTH'd2154670;
cipher_text[24] = `CIPHERTEXT_WIDTH'd15551241;
cipher_text[25] = `CIPHERTEXT_WIDTH'd6689882;
cipher_text[26] = `CIPHERTEXT_WIDTH'd12645092;
cipher_text[27] = `CIPHERTEXT_WIDTH'd13816089;
cipher_text[28] = `CIPHERTEXT_WIDTH'd4929324;
cipher_text[29] = `CIPHERTEXT_WIDTH'd1145294;
cipher_text[30] = `CIPHERTEXT_WIDTH'd14680573;
cipher_text[31] = `CIPHERTEXT_WIDTH'd4535311;
cipher_text[32] = `CIPHERTEXT_WIDTH'd9609303;
cipher_text[33] = `CIPHERTEXT_WIDTH'd2591983;
cipher_text[34] = `CIPHERTEXT_WIDTH'd10666215;
cipher_text[35] = `CIPHERTEXT_WIDTH'd14514242;
cipher_text[36] = `CIPHERTEXT_WIDTH'd9168062;
cipher_text[37] = `CIPHERTEXT_WIDTH'd1401537;
cipher_text[38] = `CIPHERTEXT_WIDTH'd6449070;
cipher_text[39] = `CIPHERTEXT_WIDTH'd7296685;
cipher_text[40] = `CIPHERTEXT_WIDTH'd13791608;
cipher_text[41] = `CIPHERTEXT_WIDTH'd15322840;
cipher_text[42] = `CIPHERTEXT_WIDTH'd16613628;
cipher_text[43] = `CIPHERTEXT_WIDTH'd3542501;
cipher_text[44] = `CIPHERTEXT_WIDTH'd16570359;
cipher_text[45] = `CIPHERTEXT_WIDTH'd3308058;
cipher_text[46] = `CIPHERTEXT_WIDTH'd514801;
cipher_text[47] = `CIPHERTEXT_WIDTH'd15000315;
cipher_text[48] = `CIPHERTEXT_WIDTH'd12333265;
cipher_text[49] = `CIPHERTEXT_WIDTH'd4159008;
cipher_text[50] = `CIPHERTEXT_WIDTH'd4305507;
cipher_text[51] = `CIPHERTEXT_WIDTH'd7327988;
cipher_text[52] = `CIPHERTEXT_WIDTH'd15549464;
cipher_text[53] = `CIPHERTEXT_WIDTH'd15108946;
cipher_text[54] = `CIPHERTEXT_WIDTH'd12000247;
cipher_text[55] = `CIPHERTEXT_WIDTH'd15442245;
cipher_text[56] = `CIPHERTEXT_WIDTH'd16679468;
cipher_text[57] = `CIPHERTEXT_WIDTH'd16482401;
cipher_text[58] = `CIPHERTEXT_WIDTH'd5373314;
cipher_text[59] = `CIPHERTEXT_WIDTH'd13765787;
cipher_text[60] = `CIPHERTEXT_WIDTH'd4560193;
cipher_text[61] = `CIPHERTEXT_WIDTH'd15439900;
cipher_text[62] = `CIPHERTEXT_WIDTH'd8684635;
cipher_text[63] = `CIPHERTEXT_WIDTH'd8109582;
cipher_text[64] = `CIPHERTEXT_WIDTH'd3369733;
cipher_text[65] = `CIPHERTEXT_WIDTH'd274628;
cipher_text[66] = `CIPHERTEXT_WIDTH'd10734831;
cipher_text[67] = `CIPHERTEXT_WIDTH'd14005783;
cipher_text[68] = `CIPHERTEXT_WIDTH'd4052706;
cipher_text[69] = `CIPHERTEXT_WIDTH'd8373224;
cipher_text[70] = `CIPHERTEXT_WIDTH'd6919308;
cipher_text[71] = `CIPHERTEXT_WIDTH'd14373598;
cipher_text[72] = `CIPHERTEXT_WIDTH'd3893790;
cipher_text[73] = `CIPHERTEXT_WIDTH'd6070219;
cipher_text[74] = `CIPHERTEXT_WIDTH'd8618683;
cipher_text[75] = `CIPHERTEXT_WIDTH'd16153353;
cipher_text[76] = `CIPHERTEXT_WIDTH'd3810814;
cipher_text[77] = `CIPHERTEXT_WIDTH'd778679;
cipher_text[78] = `CIPHERTEXT_WIDTH'd6212385;
cipher_text[79] = `CIPHERTEXT_WIDTH'd14462591;
cipher_text[80] = `CIPHERTEXT_WIDTH'd16523191;
cipher_text[81] = `CIPHERTEXT_WIDTH'd609851;
cipher_text[82] = `CIPHERTEXT_WIDTH'd4318792;
cipher_text[83] = `CIPHERTEXT_WIDTH'd7451786;
cipher_text[84] = `CIPHERTEXT_WIDTH'd4788923;
cipher_text[85] = `CIPHERTEXT_WIDTH'd13475094;
cipher_text[86] = `CIPHERTEXT_WIDTH'd2669379;
cipher_text[87] = `CIPHERTEXT_WIDTH'd6284130;
cipher_text[88] = `CIPHERTEXT_WIDTH'd6134821;
cipher_text[89] = `CIPHERTEXT_WIDTH'd4405802;
cipher_text[90] = `CIPHERTEXT_WIDTH'd14917075;
cipher_text[91] = `CIPHERTEXT_WIDTH'd5141866;
cipher_text[92] = `CIPHERTEXT_WIDTH'd16603552;
cipher_text[93] = `CIPHERTEXT_WIDTH'd4032506;
cipher_text[94] = `CIPHERTEXT_WIDTH'd13917773;
cipher_text[95] = `CIPHERTEXT_WIDTH'd7565207;
cipher_text[96] = `CIPHERTEXT_WIDTH'd14638970;
cipher_text[97] = `CIPHERTEXT_WIDTH'd5718669;
cipher_text[98] = `CIPHERTEXT_WIDTH'd9596853;
cipher_text[99] = `CIPHERTEXT_WIDTH'd10855837;
cipher_text[100] = `CIPHERTEXT_WIDTH'd16555074;
cipher_text[101] = `CIPHERTEXT_WIDTH'd8925478;
cipher_text[102] = `CIPHERTEXT_WIDTH'd4778425;
cipher_text[103] = `CIPHERTEXT_WIDTH'd7196846;
cipher_text[104] = `CIPHERTEXT_WIDTH'd6947381;
cipher_text[105] = `CIPHERTEXT_WIDTH'd3002775;
cipher_text[106] = `CIPHERTEXT_WIDTH'd15583199;
cipher_text[107] = `CIPHERTEXT_WIDTH'd10528777;
cipher_text[108] = `CIPHERTEXT_WIDTH'd15366573;
cipher_text[109] = `CIPHERTEXT_WIDTH'd1562811;
cipher_text[110] = `CIPHERTEXT_WIDTH'd3571658;
cipher_text[111] = `CIPHERTEXT_WIDTH'd15229071;
cipher_text[112] = `CIPHERTEXT_WIDTH'd2095560;
cipher_text[113] = `CIPHERTEXT_WIDTH'd238783;
cipher_text[114] = `CIPHERTEXT_WIDTH'd12003755;
cipher_text[115] = `CIPHERTEXT_WIDTH'd14996112;
cipher_text[116] = `CIPHERTEXT_WIDTH'd533395;
cipher_text[117] = `CIPHERTEXT_WIDTH'd2476013;
cipher_text[118] = `CIPHERTEXT_WIDTH'd14163690;
cipher_text[119] = `CIPHERTEXT_WIDTH'd11684021;
cipher_text[120] = `CIPHERTEXT_WIDTH'd1001177;
cipher_text[121] = `CIPHERTEXT_WIDTH'd8470014;
cipher_text[122] = `CIPHERTEXT_WIDTH'd15896918;
cipher_text[123] = `CIPHERTEXT_WIDTH'd7559099;
cipher_text[124] = `CIPHERTEXT_WIDTH'd6779456;
cipher_text[125] = `CIPHERTEXT_WIDTH'd14544966;
cipher_text[126] = `CIPHERTEXT_WIDTH'd1600598;
cipher_text[127] = `CIPHERTEXT_WIDTH'd3813055;
cipher_text[128] = `CIPHERTEXT_WIDTH'd10802891;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 15;
cipher_text[0] = `CIPHERTEXT_WIDTH'd1916185;
cipher_text[1] = `CIPHERTEXT_WIDTH'd14037304;
cipher_text[2] = `CIPHERTEXT_WIDTH'd5492599;
cipher_text[3] = `CIPHERTEXT_WIDTH'd8098517;
cipher_text[4] = `CIPHERTEXT_WIDTH'd9211629;
cipher_text[5] = `CIPHERTEXT_WIDTH'd4664444;
cipher_text[6] = `CIPHERTEXT_WIDTH'd12072964;
cipher_text[7] = `CIPHERTEXT_WIDTH'd3385920;
cipher_text[8] = `CIPHERTEXT_WIDTH'd10055909;
cipher_text[9] = `CIPHERTEXT_WIDTH'd14632308;
cipher_text[10] = `CIPHERTEXT_WIDTH'd16711426;
cipher_text[11] = `CIPHERTEXT_WIDTH'd13798066;
cipher_text[12] = `CIPHERTEXT_WIDTH'd8479331;
cipher_text[13] = `CIPHERTEXT_WIDTH'd5048564;
cipher_text[14] = `CIPHERTEXT_WIDTH'd7524530;
cipher_text[15] = `CIPHERTEXT_WIDTH'd5645162;
cipher_text[16] = `CIPHERTEXT_WIDTH'd6318171;
cipher_text[17] = `CIPHERTEXT_WIDTH'd15659322;
cipher_text[18] = `CIPHERTEXT_WIDTH'd14674779;
cipher_text[19] = `CIPHERTEXT_WIDTH'd13033132;
cipher_text[20] = `CIPHERTEXT_WIDTH'd3364891;
cipher_text[21] = `CIPHERTEXT_WIDTH'd80775;
cipher_text[22] = `CIPHERTEXT_WIDTH'd12530375;
cipher_text[23] = `CIPHERTEXT_WIDTH'd5753977;
cipher_text[24] = `CIPHERTEXT_WIDTH'd7121088;
cipher_text[25] = `CIPHERTEXT_WIDTH'd6809714;
cipher_text[26] = `CIPHERTEXT_WIDTH'd987495;
cipher_text[27] = `CIPHERTEXT_WIDTH'd13642754;
cipher_text[28] = `CIPHERTEXT_WIDTH'd2866003;
cipher_text[29] = `CIPHERTEXT_WIDTH'd3701046;
cipher_text[30] = `CIPHERTEXT_WIDTH'd14523024;
cipher_text[31] = `CIPHERTEXT_WIDTH'd2462693;
cipher_text[32] = `CIPHERTEXT_WIDTH'd9123246;
cipher_text[33] = `CIPHERTEXT_WIDTH'd8935775;
cipher_text[34] = `CIPHERTEXT_WIDTH'd4934046;
cipher_text[35] = `CIPHERTEXT_WIDTH'd14487079;
cipher_text[36] = `CIPHERTEXT_WIDTH'd7189077;
cipher_text[37] = `CIPHERTEXT_WIDTH'd6059525;
cipher_text[38] = `CIPHERTEXT_WIDTH'd14332303;
cipher_text[39] = `CIPHERTEXT_WIDTH'd15540514;
cipher_text[40] = `CIPHERTEXT_WIDTH'd12792818;
cipher_text[41] = `CIPHERTEXT_WIDTH'd3547506;
cipher_text[42] = `CIPHERTEXT_WIDTH'd5448511;
cipher_text[43] = `CIPHERTEXT_WIDTH'd8496757;
cipher_text[44] = `CIPHERTEXT_WIDTH'd7178443;
cipher_text[45] = `CIPHERTEXT_WIDTH'd2789084;
cipher_text[46] = `CIPHERTEXT_WIDTH'd13380664;
cipher_text[47] = `CIPHERTEXT_WIDTH'd3751940;
cipher_text[48] = `CIPHERTEXT_WIDTH'd16139407;
cipher_text[49] = `CIPHERTEXT_WIDTH'd12482174;
cipher_text[50] = `CIPHERTEXT_WIDTH'd5831029;
cipher_text[51] = `CIPHERTEXT_WIDTH'd3618433;
cipher_text[52] = `CIPHERTEXT_WIDTH'd14723263;
cipher_text[53] = `CIPHERTEXT_WIDTH'd6645795;
cipher_text[54] = `CIPHERTEXT_WIDTH'd8177999;
cipher_text[55] = `CIPHERTEXT_WIDTH'd4299771;
cipher_text[56] = `CIPHERTEXT_WIDTH'd1749359;
cipher_text[57] = `CIPHERTEXT_WIDTH'd16134934;
cipher_text[58] = `CIPHERTEXT_WIDTH'd1987703;
cipher_text[59] = `CIPHERTEXT_WIDTH'd4301910;
cipher_text[60] = `CIPHERTEXT_WIDTH'd6546168;
cipher_text[61] = `CIPHERTEXT_WIDTH'd10588733;
cipher_text[62] = `CIPHERTEXT_WIDTH'd10310741;
cipher_text[63] = `CIPHERTEXT_WIDTH'd7854682;
cipher_text[64] = `CIPHERTEXT_WIDTH'd1191273;
cipher_text[65] = `CIPHERTEXT_WIDTH'd11318330;
cipher_text[66] = `CIPHERTEXT_WIDTH'd12764468;
cipher_text[67] = `CIPHERTEXT_WIDTH'd701312;
cipher_text[68] = `CIPHERTEXT_WIDTH'd6090534;
cipher_text[69] = `CIPHERTEXT_WIDTH'd7414386;
cipher_text[70] = `CIPHERTEXT_WIDTH'd10283505;
cipher_text[71] = `CIPHERTEXT_WIDTH'd6455270;
cipher_text[72] = `CIPHERTEXT_WIDTH'd11922700;
cipher_text[73] = `CIPHERTEXT_WIDTH'd10891213;
cipher_text[74] = `CIPHERTEXT_WIDTH'd7771563;
cipher_text[75] = `CIPHERTEXT_WIDTH'd7023213;
cipher_text[76] = `CIPHERTEXT_WIDTH'd1598911;
cipher_text[77] = `CIPHERTEXT_WIDTH'd9460993;
cipher_text[78] = `CIPHERTEXT_WIDTH'd4027050;
cipher_text[79] = `CIPHERTEXT_WIDTH'd10994264;
cipher_text[80] = `CIPHERTEXT_WIDTH'd9338638;
cipher_text[81] = `CIPHERTEXT_WIDTH'd7336580;
cipher_text[82] = `CIPHERTEXT_WIDTH'd3985912;
cipher_text[83] = `CIPHERTEXT_WIDTH'd8539709;
cipher_text[84] = `CIPHERTEXT_WIDTH'd13421609;
cipher_text[85] = `CIPHERTEXT_WIDTH'd12159137;
cipher_text[86] = `CIPHERTEXT_WIDTH'd8654774;
cipher_text[87] = `CIPHERTEXT_WIDTH'd9054303;
cipher_text[88] = `CIPHERTEXT_WIDTH'd7624577;
cipher_text[89] = `CIPHERTEXT_WIDTH'd10015567;
cipher_text[90] = `CIPHERTEXT_WIDTH'd7324479;
cipher_text[91] = `CIPHERTEXT_WIDTH'd3707980;
cipher_text[92] = `CIPHERTEXT_WIDTH'd8833015;
cipher_text[93] = `CIPHERTEXT_WIDTH'd3176825;
cipher_text[94] = `CIPHERTEXT_WIDTH'd8485195;
cipher_text[95] = `CIPHERTEXT_WIDTH'd1018905;
cipher_text[96] = `CIPHERTEXT_WIDTH'd10338201;
cipher_text[97] = `CIPHERTEXT_WIDTH'd4926636;
cipher_text[98] = `CIPHERTEXT_WIDTH'd10952262;
cipher_text[99] = `CIPHERTEXT_WIDTH'd15475261;
cipher_text[100] = `CIPHERTEXT_WIDTH'd3612605;
cipher_text[101] = `CIPHERTEXT_WIDTH'd9396492;
cipher_text[102] = `CIPHERTEXT_WIDTH'd11620575;
cipher_text[103] = `CIPHERTEXT_WIDTH'd15426885;
cipher_text[104] = `CIPHERTEXT_WIDTH'd4346291;
cipher_text[105] = `CIPHERTEXT_WIDTH'd13586153;
cipher_text[106] = `CIPHERTEXT_WIDTH'd1691178;
cipher_text[107] = `CIPHERTEXT_WIDTH'd3936638;
cipher_text[108] = `CIPHERTEXT_WIDTH'd2697854;
cipher_text[109] = `CIPHERTEXT_WIDTH'd3306169;
cipher_text[110] = `CIPHERTEXT_WIDTH'd2616603;
cipher_text[111] = `CIPHERTEXT_WIDTH'd9662538;
cipher_text[112] = `CIPHERTEXT_WIDTH'd4818131;
cipher_text[113] = `CIPHERTEXT_WIDTH'd14926139;
cipher_text[114] = `CIPHERTEXT_WIDTH'd14604875;
cipher_text[115] = `CIPHERTEXT_WIDTH'd8359855;
cipher_text[116] = `CIPHERTEXT_WIDTH'd2169596;
cipher_text[117] = `CIPHERTEXT_WIDTH'd7252421;
cipher_text[118] = `CIPHERTEXT_WIDTH'd11526575;
cipher_text[119] = `CIPHERTEXT_WIDTH'd5737435;
cipher_text[120] = `CIPHERTEXT_WIDTH'd6135970;
cipher_text[121] = `CIPHERTEXT_WIDTH'd7108172;
cipher_text[122] = `CIPHERTEXT_WIDTH'd8286803;
cipher_text[123] = `CIPHERTEXT_WIDTH'd12297170;
cipher_text[124] = `CIPHERTEXT_WIDTH'd16613524;
cipher_text[125] = `CIPHERTEXT_WIDTH'd5282496;
cipher_text[126] = `CIPHERTEXT_WIDTH'd14876498;
cipher_text[127] = `CIPHERTEXT_WIDTH'd6148411;
cipher_text[128] = `CIPHERTEXT_WIDTH'd12903611;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 16;
cipher_text[0] = `CIPHERTEXT_WIDTH'd6740382;
cipher_text[1] = `CIPHERTEXT_WIDTH'd11454476;
cipher_text[2] = `CIPHERTEXT_WIDTH'd15994939;
cipher_text[3] = `CIPHERTEXT_WIDTH'd13186421;
cipher_text[4] = `CIPHERTEXT_WIDTH'd833345;
cipher_text[5] = `CIPHERTEXT_WIDTH'd12587166;
cipher_text[6] = `CIPHERTEXT_WIDTH'd12186664;
cipher_text[7] = `CIPHERTEXT_WIDTH'd4272644;
cipher_text[8] = `CIPHERTEXT_WIDTH'd14851637;
cipher_text[9] = `CIPHERTEXT_WIDTH'd7711499;
cipher_text[10] = `CIPHERTEXT_WIDTH'd15066095;
cipher_text[11] = `CIPHERTEXT_WIDTH'd13166166;
cipher_text[12] = `CIPHERTEXT_WIDTH'd9924474;
cipher_text[13] = `CIPHERTEXT_WIDTH'd13537632;
cipher_text[14] = `CIPHERTEXT_WIDTH'd726840;
cipher_text[15] = `CIPHERTEXT_WIDTH'd5510198;
cipher_text[16] = `CIPHERTEXT_WIDTH'd2527303;
cipher_text[17] = `CIPHERTEXT_WIDTH'd7383275;
cipher_text[18] = `CIPHERTEXT_WIDTH'd6251803;
cipher_text[19] = `CIPHERTEXT_WIDTH'd7617642;
cipher_text[20] = `CIPHERTEXT_WIDTH'd15512170;
cipher_text[21] = `CIPHERTEXT_WIDTH'd4334162;
cipher_text[22] = `CIPHERTEXT_WIDTH'd15194526;
cipher_text[23] = `CIPHERTEXT_WIDTH'd2824819;
cipher_text[24] = `CIPHERTEXT_WIDTH'd13252937;
cipher_text[25] = `CIPHERTEXT_WIDTH'd5038348;
cipher_text[26] = `CIPHERTEXT_WIDTH'd5980320;
cipher_text[27] = `CIPHERTEXT_WIDTH'd8147037;
cipher_text[28] = `CIPHERTEXT_WIDTH'd10737504;
cipher_text[29] = `CIPHERTEXT_WIDTH'd12077212;
cipher_text[30] = `CIPHERTEXT_WIDTH'd11710752;
cipher_text[31] = `CIPHERTEXT_WIDTH'd14876654;
cipher_text[32] = `CIPHERTEXT_WIDTH'd12111304;
cipher_text[33] = `CIPHERTEXT_WIDTH'd9700781;
cipher_text[34] = `CIPHERTEXT_WIDTH'd8191941;
cipher_text[35] = `CIPHERTEXT_WIDTH'd14818496;
cipher_text[36] = `CIPHERTEXT_WIDTH'd11288573;
cipher_text[37] = `CIPHERTEXT_WIDTH'd683459;
cipher_text[38] = `CIPHERTEXT_WIDTH'd1600297;
cipher_text[39] = `CIPHERTEXT_WIDTH'd6059482;
cipher_text[40] = `CIPHERTEXT_WIDTH'd12699294;
cipher_text[41] = `CIPHERTEXT_WIDTH'd6957344;
cipher_text[42] = `CIPHERTEXT_WIDTH'd2532348;
cipher_text[43] = `CIPHERTEXT_WIDTH'd9394687;
cipher_text[44] = `CIPHERTEXT_WIDTH'd5912644;
cipher_text[45] = `CIPHERTEXT_WIDTH'd8874252;
cipher_text[46] = `CIPHERTEXT_WIDTH'd5205498;
cipher_text[47] = `CIPHERTEXT_WIDTH'd7212495;
cipher_text[48] = `CIPHERTEXT_WIDTH'd14232532;
cipher_text[49] = `CIPHERTEXT_WIDTH'd1173428;
cipher_text[50] = `CIPHERTEXT_WIDTH'd2239125;
cipher_text[51] = `CIPHERTEXT_WIDTH'd4115097;
cipher_text[52] = `CIPHERTEXT_WIDTH'd14625756;
cipher_text[53] = `CIPHERTEXT_WIDTH'd12426897;
cipher_text[54] = `CIPHERTEXT_WIDTH'd11163906;
cipher_text[55] = `CIPHERTEXT_WIDTH'd11886627;
cipher_text[56] = `CIPHERTEXT_WIDTH'd7544113;
cipher_text[57] = `CIPHERTEXT_WIDTH'd5464832;
cipher_text[58] = `CIPHERTEXT_WIDTH'd2659059;
cipher_text[59] = `CIPHERTEXT_WIDTH'd8996035;
cipher_text[60] = `CIPHERTEXT_WIDTH'd5891045;
cipher_text[61] = `CIPHERTEXT_WIDTH'd13819823;
cipher_text[62] = `CIPHERTEXT_WIDTH'd15158470;
cipher_text[63] = `CIPHERTEXT_WIDTH'd11432857;
cipher_text[64] = `CIPHERTEXT_WIDTH'd12143618;
cipher_text[65] = `CIPHERTEXT_WIDTH'd6145916;
cipher_text[66] = `CIPHERTEXT_WIDTH'd358229;
cipher_text[67] = `CIPHERTEXT_WIDTH'd11045436;
cipher_text[68] = `CIPHERTEXT_WIDTH'd10759436;
cipher_text[69] = `CIPHERTEXT_WIDTH'd2910223;
cipher_text[70] = `CIPHERTEXT_WIDTH'd9701533;
cipher_text[71] = `CIPHERTEXT_WIDTH'd8256263;
cipher_text[72] = `CIPHERTEXT_WIDTH'd14956848;
cipher_text[73] = `CIPHERTEXT_WIDTH'd7443883;
cipher_text[74] = `CIPHERTEXT_WIDTH'd3806369;
cipher_text[75] = `CIPHERTEXT_WIDTH'd9259025;
cipher_text[76] = `CIPHERTEXT_WIDTH'd9710780;
cipher_text[77] = `CIPHERTEXT_WIDTH'd4107256;
cipher_text[78] = `CIPHERTEXT_WIDTH'd4315089;
cipher_text[79] = `CIPHERTEXT_WIDTH'd4752974;
cipher_text[80] = `CIPHERTEXT_WIDTH'd10194887;
cipher_text[81] = `CIPHERTEXT_WIDTH'd1498350;
cipher_text[82] = `CIPHERTEXT_WIDTH'd4946542;
cipher_text[83] = `CIPHERTEXT_WIDTH'd11949369;
cipher_text[84] = `CIPHERTEXT_WIDTH'd9150050;
cipher_text[85] = `CIPHERTEXT_WIDTH'd1141254;
cipher_text[86] = `CIPHERTEXT_WIDTH'd16650081;
cipher_text[87] = `CIPHERTEXT_WIDTH'd14746180;
cipher_text[88] = `CIPHERTEXT_WIDTH'd7624205;
cipher_text[89] = `CIPHERTEXT_WIDTH'd12776417;
cipher_text[90] = `CIPHERTEXT_WIDTH'd8156730;
cipher_text[91] = `CIPHERTEXT_WIDTH'd12875325;
cipher_text[92] = `CIPHERTEXT_WIDTH'd10479177;
cipher_text[93] = `CIPHERTEXT_WIDTH'd506575;
cipher_text[94] = `CIPHERTEXT_WIDTH'd355872;
cipher_text[95] = `CIPHERTEXT_WIDTH'd9308352;
cipher_text[96] = `CIPHERTEXT_WIDTH'd10437012;
cipher_text[97] = `CIPHERTEXT_WIDTH'd13137843;
cipher_text[98] = `CIPHERTEXT_WIDTH'd15820546;
cipher_text[99] = `CIPHERTEXT_WIDTH'd7125876;
cipher_text[100] = `CIPHERTEXT_WIDTH'd13799927;
cipher_text[101] = `CIPHERTEXT_WIDTH'd7099230;
cipher_text[102] = `CIPHERTEXT_WIDTH'd3300204;
cipher_text[103] = `CIPHERTEXT_WIDTH'd14516236;
cipher_text[104] = `CIPHERTEXT_WIDTH'd4501153;
cipher_text[105] = `CIPHERTEXT_WIDTH'd4015289;
cipher_text[106] = `CIPHERTEXT_WIDTH'd13952549;
cipher_text[107] = `CIPHERTEXT_WIDTH'd9927778;
cipher_text[108] = `CIPHERTEXT_WIDTH'd9002207;
cipher_text[109] = `CIPHERTEXT_WIDTH'd10137761;
cipher_text[110] = `CIPHERTEXT_WIDTH'd4896098;
cipher_text[111] = `CIPHERTEXT_WIDTH'd10943900;
cipher_text[112] = `CIPHERTEXT_WIDTH'd1291863;
cipher_text[113] = `CIPHERTEXT_WIDTH'd9124630;
cipher_text[114] = `CIPHERTEXT_WIDTH'd8345200;
cipher_text[115] = `CIPHERTEXT_WIDTH'd2794024;
cipher_text[116] = `CIPHERTEXT_WIDTH'd6672731;
cipher_text[117] = `CIPHERTEXT_WIDTH'd12353266;
cipher_text[118] = `CIPHERTEXT_WIDTH'd5903931;
cipher_text[119] = `CIPHERTEXT_WIDTH'd15093584;
cipher_text[120] = `CIPHERTEXT_WIDTH'd16473593;
cipher_text[121] = `CIPHERTEXT_WIDTH'd15467566;
cipher_text[122] = `CIPHERTEXT_WIDTH'd10207974;
cipher_text[123] = `CIPHERTEXT_WIDTH'd2177965;
cipher_text[124] = `CIPHERTEXT_WIDTH'd11495541;
cipher_text[125] = `CIPHERTEXT_WIDTH'd10420518;
cipher_text[126] = `CIPHERTEXT_WIDTH'd14075003;
cipher_text[127] = `CIPHERTEXT_WIDTH'd15709510;
cipher_text[128] = `CIPHERTEXT_WIDTH'd2012567;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 17;
cipher_text[0] = `CIPHERTEXT_WIDTH'd11791974;
cipher_text[1] = `CIPHERTEXT_WIDTH'd12574582;
cipher_text[2] = `CIPHERTEXT_WIDTH'd15845326;
cipher_text[3] = `CIPHERTEXT_WIDTH'd964047;
cipher_text[4] = `CIPHERTEXT_WIDTH'd5563256;
cipher_text[5] = `CIPHERTEXT_WIDTH'd1895598;
cipher_text[6] = `CIPHERTEXT_WIDTH'd4132619;
cipher_text[7] = `CIPHERTEXT_WIDTH'd14985544;
cipher_text[8] = `CIPHERTEXT_WIDTH'd2786701;
cipher_text[9] = `CIPHERTEXT_WIDTH'd10261361;
cipher_text[10] = `CIPHERTEXT_WIDTH'd1501044;
cipher_text[11] = `CIPHERTEXT_WIDTH'd4957753;
cipher_text[12] = `CIPHERTEXT_WIDTH'd5826377;
cipher_text[13] = `CIPHERTEXT_WIDTH'd6974074;
cipher_text[14] = `CIPHERTEXT_WIDTH'd3071895;
cipher_text[15] = `CIPHERTEXT_WIDTH'd2587358;
cipher_text[16] = `CIPHERTEXT_WIDTH'd8721475;
cipher_text[17] = `CIPHERTEXT_WIDTH'd7952563;
cipher_text[18] = `CIPHERTEXT_WIDTH'd16179416;
cipher_text[19] = `CIPHERTEXT_WIDTH'd4057637;
cipher_text[20] = `CIPHERTEXT_WIDTH'd15851381;
cipher_text[21] = `CIPHERTEXT_WIDTH'd4017967;
cipher_text[22] = `CIPHERTEXT_WIDTH'd8156495;
cipher_text[23] = `CIPHERTEXT_WIDTH'd10942483;
cipher_text[24] = `CIPHERTEXT_WIDTH'd3693293;
cipher_text[25] = `CIPHERTEXT_WIDTH'd51506;
cipher_text[26] = `CIPHERTEXT_WIDTH'd4449108;
cipher_text[27] = `CIPHERTEXT_WIDTH'd2589540;
cipher_text[28] = `CIPHERTEXT_WIDTH'd16396223;
cipher_text[29] = `CIPHERTEXT_WIDTH'd9340085;
cipher_text[30] = `CIPHERTEXT_WIDTH'd6877483;
cipher_text[31] = `CIPHERTEXT_WIDTH'd15310541;
cipher_text[32] = `CIPHERTEXT_WIDTH'd15089184;
cipher_text[33] = `CIPHERTEXT_WIDTH'd3555643;
cipher_text[34] = `CIPHERTEXT_WIDTH'd13634453;
cipher_text[35] = `CIPHERTEXT_WIDTH'd13093579;
cipher_text[36] = `CIPHERTEXT_WIDTH'd10564454;
cipher_text[37] = `CIPHERTEXT_WIDTH'd13436210;
cipher_text[38] = `CIPHERTEXT_WIDTH'd3049709;
cipher_text[39] = `CIPHERTEXT_WIDTH'd6587727;
cipher_text[40] = `CIPHERTEXT_WIDTH'd5724292;
cipher_text[41] = `CIPHERTEXT_WIDTH'd10179359;
cipher_text[42] = `CIPHERTEXT_WIDTH'd9295467;
cipher_text[43] = `CIPHERTEXT_WIDTH'd10453839;
cipher_text[44] = `CIPHERTEXT_WIDTH'd11297387;
cipher_text[45] = `CIPHERTEXT_WIDTH'd10851396;
cipher_text[46] = `CIPHERTEXT_WIDTH'd2003606;
cipher_text[47] = `CIPHERTEXT_WIDTH'd4296511;
cipher_text[48] = `CIPHERTEXT_WIDTH'd8166705;
cipher_text[49] = `CIPHERTEXT_WIDTH'd8429486;
cipher_text[50] = `CIPHERTEXT_WIDTH'd9639575;
cipher_text[51] = `CIPHERTEXT_WIDTH'd11364727;
cipher_text[52] = `CIPHERTEXT_WIDTH'd7116187;
cipher_text[53] = `CIPHERTEXT_WIDTH'd14079466;
cipher_text[54] = `CIPHERTEXT_WIDTH'd4873492;
cipher_text[55] = `CIPHERTEXT_WIDTH'd10986752;
cipher_text[56] = `CIPHERTEXT_WIDTH'd10078259;
cipher_text[57] = `CIPHERTEXT_WIDTH'd9560192;
cipher_text[58] = `CIPHERTEXT_WIDTH'd16538509;
cipher_text[59] = `CIPHERTEXT_WIDTH'd6297136;
cipher_text[60] = `CIPHERTEXT_WIDTH'd1291374;
cipher_text[61] = `CIPHERTEXT_WIDTH'd7485099;
cipher_text[62] = `CIPHERTEXT_WIDTH'd9898122;
cipher_text[63] = `CIPHERTEXT_WIDTH'd2943674;
cipher_text[64] = `CIPHERTEXT_WIDTH'd7121053;
cipher_text[65] = `CIPHERTEXT_WIDTH'd7754211;
cipher_text[66] = `CIPHERTEXT_WIDTH'd8188077;
cipher_text[67] = `CIPHERTEXT_WIDTH'd7559885;
cipher_text[68] = `CIPHERTEXT_WIDTH'd5736228;
cipher_text[69] = `CIPHERTEXT_WIDTH'd14794062;
cipher_text[70] = `CIPHERTEXT_WIDTH'd1481975;
cipher_text[71] = `CIPHERTEXT_WIDTH'd6765925;
cipher_text[72] = `CIPHERTEXT_WIDTH'd7319599;
cipher_text[73] = `CIPHERTEXT_WIDTH'd5377066;
cipher_text[74] = `CIPHERTEXT_WIDTH'd15766894;
cipher_text[75] = `CIPHERTEXT_WIDTH'd14781949;
cipher_text[76] = `CIPHERTEXT_WIDTH'd9650335;
cipher_text[77] = `CIPHERTEXT_WIDTH'd15646396;
cipher_text[78] = `CIPHERTEXT_WIDTH'd12849055;
cipher_text[79] = `CIPHERTEXT_WIDTH'd1718509;
cipher_text[80] = `CIPHERTEXT_WIDTH'd8235750;
cipher_text[81] = `CIPHERTEXT_WIDTH'd7933798;
cipher_text[82] = `CIPHERTEXT_WIDTH'd10288977;
cipher_text[83] = `CIPHERTEXT_WIDTH'd1646187;
cipher_text[84] = `CIPHERTEXT_WIDTH'd13912463;
cipher_text[85] = `CIPHERTEXT_WIDTH'd6932218;
cipher_text[86] = `CIPHERTEXT_WIDTH'd13685012;
cipher_text[87] = `CIPHERTEXT_WIDTH'd9828917;
cipher_text[88] = `CIPHERTEXT_WIDTH'd7611728;
cipher_text[89] = `CIPHERTEXT_WIDTH'd3446589;
cipher_text[90] = `CIPHERTEXT_WIDTH'd14209984;
cipher_text[91] = `CIPHERTEXT_WIDTH'd11563584;
cipher_text[92] = `CIPHERTEXT_WIDTH'd2614938;
cipher_text[93] = `CIPHERTEXT_WIDTH'd1269267;
cipher_text[94] = `CIPHERTEXT_WIDTH'd9647835;
cipher_text[95] = `CIPHERTEXT_WIDTH'd12796316;
cipher_text[96] = `CIPHERTEXT_WIDTH'd8676053;
cipher_text[97] = `CIPHERTEXT_WIDTH'd12544679;
cipher_text[98] = `CIPHERTEXT_WIDTH'd13871651;
cipher_text[99] = `CIPHERTEXT_WIDTH'd11575559;
cipher_text[100] = `CIPHERTEXT_WIDTH'd13036497;
cipher_text[101] = `CIPHERTEXT_WIDTH'd11445411;
cipher_text[102] = `CIPHERTEXT_WIDTH'd1718478;
cipher_text[103] = `CIPHERTEXT_WIDTH'd6654814;
cipher_text[104] = `CIPHERTEXT_WIDTH'd5540526;
cipher_text[105] = `CIPHERTEXT_WIDTH'd5234140;
cipher_text[106] = `CIPHERTEXT_WIDTH'd16116553;
cipher_text[107] = `CIPHERTEXT_WIDTH'd5878194;
cipher_text[108] = `CIPHERTEXT_WIDTH'd6346231;
cipher_text[109] = `CIPHERTEXT_WIDTH'd3264701;
cipher_text[110] = `CIPHERTEXT_WIDTH'd16495370;
cipher_text[111] = `CIPHERTEXT_WIDTH'd6338838;
cipher_text[112] = `CIPHERTEXT_WIDTH'd14583340;
cipher_text[113] = `CIPHERTEXT_WIDTH'd11221496;
cipher_text[114] = `CIPHERTEXT_WIDTH'd7122530;
cipher_text[115] = `CIPHERTEXT_WIDTH'd16577611;
cipher_text[116] = `CIPHERTEXT_WIDTH'd3978460;
cipher_text[117] = `CIPHERTEXT_WIDTH'd11475869;
cipher_text[118] = `CIPHERTEXT_WIDTH'd13538896;
cipher_text[119] = `CIPHERTEXT_WIDTH'd11297485;
cipher_text[120] = `CIPHERTEXT_WIDTH'd6475178;
cipher_text[121] = `CIPHERTEXT_WIDTH'd9053314;
cipher_text[122] = `CIPHERTEXT_WIDTH'd6483931;
cipher_text[123] = `CIPHERTEXT_WIDTH'd3935474;
cipher_text[124] = `CIPHERTEXT_WIDTH'd5509099;
cipher_text[125] = `CIPHERTEXT_WIDTH'd3434395;
cipher_text[126] = `CIPHERTEXT_WIDTH'd12501500;
cipher_text[127] = `CIPHERTEXT_WIDTH'd6592800;
cipher_text[128] = `CIPHERTEXT_WIDTH'd3496852;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 18;
cipher_text[0] = `CIPHERTEXT_WIDTH'd12998312;
cipher_text[1] = `CIPHERTEXT_WIDTH'd15449472;
cipher_text[2] = `CIPHERTEXT_WIDTH'd11517080;
cipher_text[3] = `CIPHERTEXT_WIDTH'd12444511;
cipher_text[4] = `CIPHERTEXT_WIDTH'd9409984;
cipher_text[5] = `CIPHERTEXT_WIDTH'd10681398;
cipher_text[6] = `CIPHERTEXT_WIDTH'd12268936;
cipher_text[7] = `CIPHERTEXT_WIDTH'd4140795;
cipher_text[8] = `CIPHERTEXT_WIDTH'd15192486;
cipher_text[9] = `CIPHERTEXT_WIDTH'd5192069;
cipher_text[10] = `CIPHERTEXT_WIDTH'd12705297;
cipher_text[11] = `CIPHERTEXT_WIDTH'd8876974;
cipher_text[12] = `CIPHERTEXT_WIDTH'd1196071;
cipher_text[13] = `CIPHERTEXT_WIDTH'd13210266;
cipher_text[14] = `CIPHERTEXT_WIDTH'd10201009;
cipher_text[15] = `CIPHERTEXT_WIDTH'd469817;
cipher_text[16] = `CIPHERTEXT_WIDTH'd179704;
cipher_text[17] = `CIPHERTEXT_WIDTH'd9025116;
cipher_text[18] = `CIPHERTEXT_WIDTH'd8472360;
cipher_text[19] = `CIPHERTEXT_WIDTH'd13041373;
cipher_text[20] = `CIPHERTEXT_WIDTH'd2728142;
cipher_text[21] = `CIPHERTEXT_WIDTH'd11292056;
cipher_text[22] = `CIPHERTEXT_WIDTH'd2966928;
cipher_text[23] = `CIPHERTEXT_WIDTH'd12739379;
cipher_text[24] = `CIPHERTEXT_WIDTH'd8773814;
cipher_text[25] = `CIPHERTEXT_WIDTH'd16701141;
cipher_text[26] = `CIPHERTEXT_WIDTH'd2258654;
cipher_text[27] = `CIPHERTEXT_WIDTH'd5715809;
cipher_text[28] = `CIPHERTEXT_WIDTH'd2916291;
cipher_text[29] = `CIPHERTEXT_WIDTH'd2124613;
cipher_text[30] = `CIPHERTEXT_WIDTH'd4982300;
cipher_text[31] = `CIPHERTEXT_WIDTH'd664301;
cipher_text[32] = `CIPHERTEXT_WIDTH'd6337429;
cipher_text[33] = `CIPHERTEXT_WIDTH'd7128950;
cipher_text[34] = `CIPHERTEXT_WIDTH'd11667764;
cipher_text[35] = `CIPHERTEXT_WIDTH'd6401445;
cipher_text[36] = `CIPHERTEXT_WIDTH'd1610229;
cipher_text[37] = `CIPHERTEXT_WIDTH'd12259123;
cipher_text[38] = `CIPHERTEXT_WIDTH'd8112331;
cipher_text[39] = `CIPHERTEXT_WIDTH'd13882927;
cipher_text[40] = `CIPHERTEXT_WIDTH'd13346750;
cipher_text[41] = `CIPHERTEXT_WIDTH'd4329816;
cipher_text[42] = `CIPHERTEXT_WIDTH'd1662287;
cipher_text[43] = `CIPHERTEXT_WIDTH'd8278320;
cipher_text[44] = `CIPHERTEXT_WIDTH'd4268614;
cipher_text[45] = `CIPHERTEXT_WIDTH'd7043659;
cipher_text[46] = `CIPHERTEXT_WIDTH'd12283030;
cipher_text[47] = `CIPHERTEXT_WIDTH'd9248437;
cipher_text[48] = `CIPHERTEXT_WIDTH'd16639267;
cipher_text[49] = `CIPHERTEXT_WIDTH'd10824449;
cipher_text[50] = `CIPHERTEXT_WIDTH'd2812607;
cipher_text[51] = `CIPHERTEXT_WIDTH'd12439258;
cipher_text[52] = `CIPHERTEXT_WIDTH'd11652173;
cipher_text[53] = `CIPHERTEXT_WIDTH'd3516699;
cipher_text[54] = `CIPHERTEXT_WIDTH'd11457851;
cipher_text[55] = `CIPHERTEXT_WIDTH'd10946411;
cipher_text[56] = `CIPHERTEXT_WIDTH'd13675671;
cipher_text[57] = `CIPHERTEXT_WIDTH'd11369111;
cipher_text[58] = `CIPHERTEXT_WIDTH'd9194370;
cipher_text[59] = `CIPHERTEXT_WIDTH'd1563554;
cipher_text[60] = `CIPHERTEXT_WIDTH'd3181414;
cipher_text[61] = `CIPHERTEXT_WIDTH'd3122175;
cipher_text[62] = `CIPHERTEXT_WIDTH'd9247088;
cipher_text[63] = `CIPHERTEXT_WIDTH'd9790498;
cipher_text[64] = `CIPHERTEXT_WIDTH'd11622434;
cipher_text[65] = `CIPHERTEXT_WIDTH'd184721;
cipher_text[66] = `CIPHERTEXT_WIDTH'd563770;
cipher_text[67] = `CIPHERTEXT_WIDTH'd9026903;
cipher_text[68] = `CIPHERTEXT_WIDTH'd9131599;
cipher_text[69] = `CIPHERTEXT_WIDTH'd12599614;
cipher_text[70] = `CIPHERTEXT_WIDTH'd4769220;
cipher_text[71] = `CIPHERTEXT_WIDTH'd14609107;
cipher_text[72] = `CIPHERTEXT_WIDTH'd6359811;
cipher_text[73] = `CIPHERTEXT_WIDTH'd7530440;
cipher_text[74] = `CIPHERTEXT_WIDTH'd5766019;
cipher_text[75] = `CIPHERTEXT_WIDTH'd6573746;
cipher_text[76] = `CIPHERTEXT_WIDTH'd15392671;
cipher_text[77] = `CIPHERTEXT_WIDTH'd579642;
cipher_text[78] = `CIPHERTEXT_WIDTH'd3359899;
cipher_text[79] = `CIPHERTEXT_WIDTH'd9803654;
cipher_text[80] = `CIPHERTEXT_WIDTH'd6308650;
cipher_text[81] = `CIPHERTEXT_WIDTH'd4393095;
cipher_text[82] = `CIPHERTEXT_WIDTH'd3752099;
cipher_text[83] = `CIPHERTEXT_WIDTH'd8959660;
cipher_text[84] = `CIPHERTEXT_WIDTH'd13571228;
cipher_text[85] = `CIPHERTEXT_WIDTH'd5014783;
cipher_text[86] = `CIPHERTEXT_WIDTH'd3387034;
cipher_text[87] = `CIPHERTEXT_WIDTH'd11572906;
cipher_text[88] = `CIPHERTEXT_WIDTH'd2382351;
cipher_text[89] = `CIPHERTEXT_WIDTH'd10847193;
cipher_text[90] = `CIPHERTEXT_WIDTH'd3254962;
cipher_text[91] = `CIPHERTEXT_WIDTH'd5349287;
cipher_text[92] = `CIPHERTEXT_WIDTH'd2206585;
cipher_text[93] = `CIPHERTEXT_WIDTH'd12960052;
cipher_text[94] = `CIPHERTEXT_WIDTH'd10546029;
cipher_text[95] = `CIPHERTEXT_WIDTH'd3127924;
cipher_text[96] = `CIPHERTEXT_WIDTH'd3999274;
cipher_text[97] = `CIPHERTEXT_WIDTH'd12892813;
cipher_text[98] = `CIPHERTEXT_WIDTH'd2901356;
cipher_text[99] = `CIPHERTEXT_WIDTH'd236580;
cipher_text[100] = `CIPHERTEXT_WIDTH'd8524910;
cipher_text[101] = `CIPHERTEXT_WIDTH'd3356517;
cipher_text[102] = `CIPHERTEXT_WIDTH'd15123201;
cipher_text[103] = `CIPHERTEXT_WIDTH'd15328315;
cipher_text[104] = `CIPHERTEXT_WIDTH'd9917998;
cipher_text[105] = `CIPHERTEXT_WIDTH'd16756391;
cipher_text[106] = `CIPHERTEXT_WIDTH'd1445552;
cipher_text[107] = `CIPHERTEXT_WIDTH'd4339023;
cipher_text[108] = `CIPHERTEXT_WIDTH'd10364175;
cipher_text[109] = `CIPHERTEXT_WIDTH'd2942034;
cipher_text[110] = `CIPHERTEXT_WIDTH'd14141160;
cipher_text[111] = `CIPHERTEXT_WIDTH'd13756458;
cipher_text[112] = `CIPHERTEXT_WIDTH'd4723447;
cipher_text[113] = `CIPHERTEXT_WIDTH'd282536;
cipher_text[114] = `CIPHERTEXT_WIDTH'd7485963;
cipher_text[115] = `CIPHERTEXT_WIDTH'd3509768;
cipher_text[116] = `CIPHERTEXT_WIDTH'd7311842;
cipher_text[117] = `CIPHERTEXT_WIDTH'd7506659;
cipher_text[118] = `CIPHERTEXT_WIDTH'd15234094;
cipher_text[119] = `CIPHERTEXT_WIDTH'd4422093;
cipher_text[120] = `CIPHERTEXT_WIDTH'd1990865;
cipher_text[121] = `CIPHERTEXT_WIDTH'd1926041;
cipher_text[122] = `CIPHERTEXT_WIDTH'd6017917;
cipher_text[123] = `CIPHERTEXT_WIDTH'd2099562;
cipher_text[124] = `CIPHERTEXT_WIDTH'd5300143;
cipher_text[125] = `CIPHERTEXT_WIDTH'd8481995;
cipher_text[126] = `CIPHERTEXT_WIDTH'd11072007;
cipher_text[127] = `CIPHERTEXT_WIDTH'd2522339;
cipher_text[128] = `CIPHERTEXT_WIDTH'd15482108;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 19;
cipher_text[0] = `CIPHERTEXT_WIDTH'd4845800;
cipher_text[1] = `CIPHERTEXT_WIDTH'd10137109;
cipher_text[2] = `CIPHERTEXT_WIDTH'd2695606;
cipher_text[3] = `CIPHERTEXT_WIDTH'd11407188;
cipher_text[4] = `CIPHERTEXT_WIDTH'd46829;
cipher_text[5] = `CIPHERTEXT_WIDTH'd8070364;
cipher_text[6] = `CIPHERTEXT_WIDTH'd10244017;
cipher_text[7] = `CIPHERTEXT_WIDTH'd10340600;
cipher_text[8] = `CIPHERTEXT_WIDTH'd13442189;
cipher_text[9] = `CIPHERTEXT_WIDTH'd3499979;
cipher_text[10] = `CIPHERTEXT_WIDTH'd12133638;
cipher_text[11] = `CIPHERTEXT_WIDTH'd9688863;
cipher_text[12] = `CIPHERTEXT_WIDTH'd16434982;
cipher_text[13] = `CIPHERTEXT_WIDTH'd16216072;
cipher_text[14] = `CIPHERTEXT_WIDTH'd1773703;
cipher_text[15] = `CIPHERTEXT_WIDTH'd7215927;
cipher_text[16] = `CIPHERTEXT_WIDTH'd1772700;
cipher_text[17] = `CIPHERTEXT_WIDTH'd9597553;
cipher_text[18] = `CIPHERTEXT_WIDTH'd1996882;
cipher_text[19] = `CIPHERTEXT_WIDTH'd15301889;
cipher_text[20] = `CIPHERTEXT_WIDTH'd2128301;
cipher_text[21] = `CIPHERTEXT_WIDTH'd13670176;
cipher_text[22] = `CIPHERTEXT_WIDTH'd14350518;
cipher_text[23] = `CIPHERTEXT_WIDTH'd3528218;
cipher_text[24] = `CIPHERTEXT_WIDTH'd3486150;
cipher_text[25] = `CIPHERTEXT_WIDTH'd6656777;
cipher_text[26] = `CIPHERTEXT_WIDTH'd15427328;
cipher_text[27] = `CIPHERTEXT_WIDTH'd6082516;
cipher_text[28] = `CIPHERTEXT_WIDTH'd9964838;
cipher_text[29] = `CIPHERTEXT_WIDTH'd11080009;
cipher_text[30] = `CIPHERTEXT_WIDTH'd8930973;
cipher_text[31] = `CIPHERTEXT_WIDTH'd9669073;
cipher_text[32] = `CIPHERTEXT_WIDTH'd5211531;
cipher_text[33] = `CIPHERTEXT_WIDTH'd11819953;
cipher_text[34] = `CIPHERTEXT_WIDTH'd4498660;
cipher_text[35] = `CIPHERTEXT_WIDTH'd3501135;
cipher_text[36] = `CIPHERTEXT_WIDTH'd9962422;
cipher_text[37] = `CIPHERTEXT_WIDTH'd15735312;
cipher_text[38] = `CIPHERTEXT_WIDTH'd6840118;
cipher_text[39] = `CIPHERTEXT_WIDTH'd9341354;
cipher_text[40] = `CIPHERTEXT_WIDTH'd14911407;
cipher_text[41] = `CIPHERTEXT_WIDTH'd12583808;
cipher_text[42] = `CIPHERTEXT_WIDTH'd15805061;
cipher_text[43] = `CIPHERTEXT_WIDTH'd4347248;
cipher_text[44] = `CIPHERTEXT_WIDTH'd8194162;
cipher_text[45] = `CIPHERTEXT_WIDTH'd6426032;
cipher_text[46] = `CIPHERTEXT_WIDTH'd12069158;
cipher_text[47] = `CIPHERTEXT_WIDTH'd9950641;
cipher_text[48] = `CIPHERTEXT_WIDTH'd10113231;
cipher_text[49] = `CIPHERTEXT_WIDTH'd10498957;
cipher_text[50] = `CIPHERTEXT_WIDTH'd9208543;
cipher_text[51] = `CIPHERTEXT_WIDTH'd8023710;
cipher_text[52] = `CIPHERTEXT_WIDTH'd3929743;
cipher_text[53] = `CIPHERTEXT_WIDTH'd8843549;
cipher_text[54] = `CIPHERTEXT_WIDTH'd5979335;
cipher_text[55] = `CIPHERTEXT_WIDTH'd14372688;
cipher_text[56] = `CIPHERTEXT_WIDTH'd15025307;
cipher_text[57] = `CIPHERTEXT_WIDTH'd8230296;
cipher_text[58] = `CIPHERTEXT_WIDTH'd14543780;
cipher_text[59] = `CIPHERTEXT_WIDTH'd11032586;
cipher_text[60] = `CIPHERTEXT_WIDTH'd10937680;
cipher_text[61] = `CIPHERTEXT_WIDTH'd6764396;
cipher_text[62] = `CIPHERTEXT_WIDTH'd16260578;
cipher_text[63] = `CIPHERTEXT_WIDTH'd3536335;
cipher_text[64] = `CIPHERTEXT_WIDTH'd8258776;
cipher_text[65] = `CIPHERTEXT_WIDTH'd1052363;
cipher_text[66] = `CIPHERTEXT_WIDTH'd9102189;
cipher_text[67] = `CIPHERTEXT_WIDTH'd1211309;
cipher_text[68] = `CIPHERTEXT_WIDTH'd16683652;
cipher_text[69] = `CIPHERTEXT_WIDTH'd6117354;
cipher_text[70] = `CIPHERTEXT_WIDTH'd1539811;
cipher_text[71] = `CIPHERTEXT_WIDTH'd10824402;
cipher_text[72] = `CIPHERTEXT_WIDTH'd16766221;
cipher_text[73] = `CIPHERTEXT_WIDTH'd7283462;
cipher_text[74] = `CIPHERTEXT_WIDTH'd751646;
cipher_text[75] = `CIPHERTEXT_WIDTH'd3552002;
cipher_text[76] = `CIPHERTEXT_WIDTH'd2771824;
cipher_text[77] = `CIPHERTEXT_WIDTH'd13527944;
cipher_text[78] = `CIPHERTEXT_WIDTH'd16546985;
cipher_text[79] = `CIPHERTEXT_WIDTH'd16159035;
cipher_text[80] = `CIPHERTEXT_WIDTH'd8808859;
cipher_text[81] = `CIPHERTEXT_WIDTH'd13410581;
cipher_text[82] = `CIPHERTEXT_WIDTH'd6365704;
cipher_text[83] = `CIPHERTEXT_WIDTH'd8047095;
cipher_text[84] = `CIPHERTEXT_WIDTH'd14039298;
cipher_text[85] = `CIPHERTEXT_WIDTH'd949480;
cipher_text[86] = `CIPHERTEXT_WIDTH'd1368845;
cipher_text[87] = `CIPHERTEXT_WIDTH'd2130158;
cipher_text[88] = `CIPHERTEXT_WIDTH'd1160911;
cipher_text[89] = `CIPHERTEXT_WIDTH'd4659846;
cipher_text[90] = `CIPHERTEXT_WIDTH'd14475388;
cipher_text[91] = `CIPHERTEXT_WIDTH'd12116895;
cipher_text[92] = `CIPHERTEXT_WIDTH'd6541674;
cipher_text[93] = `CIPHERTEXT_WIDTH'd3830961;
cipher_text[94] = `CIPHERTEXT_WIDTH'd15152711;
cipher_text[95] = `CIPHERTEXT_WIDTH'd8415592;
cipher_text[96] = `CIPHERTEXT_WIDTH'd5639941;
cipher_text[97] = `CIPHERTEXT_WIDTH'd5950518;
cipher_text[98] = `CIPHERTEXT_WIDTH'd9048473;
cipher_text[99] = `CIPHERTEXT_WIDTH'd4115428;
cipher_text[100] = `CIPHERTEXT_WIDTH'd4991140;
cipher_text[101] = `CIPHERTEXT_WIDTH'd3367424;
cipher_text[102] = `CIPHERTEXT_WIDTH'd13489124;
cipher_text[103] = `CIPHERTEXT_WIDTH'd5120078;
cipher_text[104] = `CIPHERTEXT_WIDTH'd9144755;
cipher_text[105] = `CIPHERTEXT_WIDTH'd10628997;
cipher_text[106] = `CIPHERTEXT_WIDTH'd13592271;
cipher_text[107] = `CIPHERTEXT_WIDTH'd12974657;
cipher_text[108] = `CIPHERTEXT_WIDTH'd8638924;
cipher_text[109] = `CIPHERTEXT_WIDTH'd2288127;
cipher_text[110] = `CIPHERTEXT_WIDTH'd3792347;
cipher_text[111] = `CIPHERTEXT_WIDTH'd1503296;
cipher_text[112] = `CIPHERTEXT_WIDTH'd11249028;
cipher_text[113] = `CIPHERTEXT_WIDTH'd15219408;
cipher_text[114] = `CIPHERTEXT_WIDTH'd10264808;
cipher_text[115] = `CIPHERTEXT_WIDTH'd15267351;
cipher_text[116] = `CIPHERTEXT_WIDTH'd5177229;
cipher_text[117] = `CIPHERTEXT_WIDTH'd5021351;
cipher_text[118] = `CIPHERTEXT_WIDTH'd3572224;
cipher_text[119] = `CIPHERTEXT_WIDTH'd3648844;
cipher_text[120] = `CIPHERTEXT_WIDTH'd12519482;
cipher_text[121] = `CIPHERTEXT_WIDTH'd6406128;
cipher_text[122] = `CIPHERTEXT_WIDTH'd15424865;
cipher_text[123] = `CIPHERTEXT_WIDTH'd8560814;
cipher_text[124] = `CIPHERTEXT_WIDTH'd2001914;
cipher_text[125] = `CIPHERTEXT_WIDTH'd7399192;
cipher_text[126] = `CIPHERTEXT_WIDTH'd13548390;
cipher_text[127] = `CIPHERTEXT_WIDTH'd942206;
cipher_text[128] = `CIPHERTEXT_WIDTH'd15449823;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 20;
cipher_text[0] = `CIPHERTEXT_WIDTH'd14987191;
cipher_text[1] = `CIPHERTEXT_WIDTH'd7847825;
cipher_text[2] = `CIPHERTEXT_WIDTH'd9157954;
cipher_text[3] = `CIPHERTEXT_WIDTH'd7609283;
cipher_text[4] = `CIPHERTEXT_WIDTH'd2646952;
cipher_text[5] = `CIPHERTEXT_WIDTH'd5955891;
cipher_text[6] = `CIPHERTEXT_WIDTH'd2899116;
cipher_text[7] = `CIPHERTEXT_WIDTH'd2025631;
cipher_text[8] = `CIPHERTEXT_WIDTH'd10942896;
cipher_text[9] = `CIPHERTEXT_WIDTH'd16400509;
cipher_text[10] = `CIPHERTEXT_WIDTH'd16079505;
cipher_text[11] = `CIPHERTEXT_WIDTH'd9315781;
cipher_text[12] = `CIPHERTEXT_WIDTH'd13889842;
cipher_text[13] = `CIPHERTEXT_WIDTH'd3587004;
cipher_text[14] = `CIPHERTEXT_WIDTH'd5063652;
cipher_text[15] = `CIPHERTEXT_WIDTH'd3489575;
cipher_text[16] = `CIPHERTEXT_WIDTH'd9644835;
cipher_text[17] = `CIPHERTEXT_WIDTH'd5374031;
cipher_text[18] = `CIPHERTEXT_WIDTH'd9854415;
cipher_text[19] = `CIPHERTEXT_WIDTH'd15413448;
cipher_text[20] = `CIPHERTEXT_WIDTH'd3705585;
cipher_text[21] = `CIPHERTEXT_WIDTH'd814018;
cipher_text[22] = `CIPHERTEXT_WIDTH'd969427;
cipher_text[23] = `CIPHERTEXT_WIDTH'd3213189;
cipher_text[24] = `CIPHERTEXT_WIDTH'd8917808;
cipher_text[25] = `CIPHERTEXT_WIDTH'd2980061;
cipher_text[26] = `CIPHERTEXT_WIDTH'd2813577;
cipher_text[27] = `CIPHERTEXT_WIDTH'd8922099;
cipher_text[28] = `CIPHERTEXT_WIDTH'd6395141;
cipher_text[29] = `CIPHERTEXT_WIDTH'd8013952;
cipher_text[30] = `CIPHERTEXT_WIDTH'd10308706;
cipher_text[31] = `CIPHERTEXT_WIDTH'd12475146;
cipher_text[32] = `CIPHERTEXT_WIDTH'd9860943;
cipher_text[33] = `CIPHERTEXT_WIDTH'd535682;
cipher_text[34] = `CIPHERTEXT_WIDTH'd10496232;
cipher_text[35] = `CIPHERTEXT_WIDTH'd16512827;
cipher_text[36] = `CIPHERTEXT_WIDTH'd11164406;
cipher_text[37] = `CIPHERTEXT_WIDTH'd16611918;
cipher_text[38] = `CIPHERTEXT_WIDTH'd11235677;
cipher_text[39] = `CIPHERTEXT_WIDTH'd5756409;
cipher_text[40] = `CIPHERTEXT_WIDTH'd2057963;
cipher_text[41] = `CIPHERTEXT_WIDTH'd4691026;
cipher_text[42] = `CIPHERTEXT_WIDTH'd3674596;
cipher_text[43] = `CIPHERTEXT_WIDTH'd12486899;
cipher_text[44] = `CIPHERTEXT_WIDTH'd5305949;
cipher_text[45] = `CIPHERTEXT_WIDTH'd4441545;
cipher_text[46] = `CIPHERTEXT_WIDTH'd11325042;
cipher_text[47] = `CIPHERTEXT_WIDTH'd4207756;
cipher_text[48] = `CIPHERTEXT_WIDTH'd4172474;
cipher_text[49] = `CIPHERTEXT_WIDTH'd9779088;
cipher_text[50] = `CIPHERTEXT_WIDTH'd2746486;
cipher_text[51] = `CIPHERTEXT_WIDTH'd1571054;
cipher_text[52] = `CIPHERTEXT_WIDTH'd2173248;
cipher_text[53] = `CIPHERTEXT_WIDTH'd16632711;
cipher_text[54] = `CIPHERTEXT_WIDTH'd12068534;
cipher_text[55] = `CIPHERTEXT_WIDTH'd13399633;
cipher_text[56] = `CIPHERTEXT_WIDTH'd9595049;
cipher_text[57] = `CIPHERTEXT_WIDTH'd3910893;
cipher_text[58] = `CIPHERTEXT_WIDTH'd11164182;
cipher_text[59] = `CIPHERTEXT_WIDTH'd14752696;
cipher_text[60] = `CIPHERTEXT_WIDTH'd13153351;
cipher_text[61] = `CIPHERTEXT_WIDTH'd15356412;
cipher_text[62] = `CIPHERTEXT_WIDTH'd15209667;
cipher_text[63] = `CIPHERTEXT_WIDTH'd7689852;
cipher_text[64] = `CIPHERTEXT_WIDTH'd8567970;
cipher_text[65] = `CIPHERTEXT_WIDTH'd15144009;
cipher_text[66] = `CIPHERTEXT_WIDTH'd16525730;
cipher_text[67] = `CIPHERTEXT_WIDTH'd3959286;
cipher_text[68] = `CIPHERTEXT_WIDTH'd1937426;
cipher_text[69] = `CIPHERTEXT_WIDTH'd3437296;
cipher_text[70] = `CIPHERTEXT_WIDTH'd6998306;
cipher_text[71] = `CIPHERTEXT_WIDTH'd12960003;
cipher_text[72] = `CIPHERTEXT_WIDTH'd9742024;
cipher_text[73] = `CIPHERTEXT_WIDTH'd672699;
cipher_text[74] = `CIPHERTEXT_WIDTH'd15026761;
cipher_text[75] = `CIPHERTEXT_WIDTH'd1536250;
cipher_text[76] = `CIPHERTEXT_WIDTH'd10755654;
cipher_text[77] = `CIPHERTEXT_WIDTH'd6640428;
cipher_text[78] = `CIPHERTEXT_WIDTH'd3166573;
cipher_text[79] = `CIPHERTEXT_WIDTH'd5711653;
cipher_text[80] = `CIPHERTEXT_WIDTH'd3771235;
cipher_text[81] = `CIPHERTEXT_WIDTH'd6344676;
cipher_text[82] = `CIPHERTEXT_WIDTH'd6446512;
cipher_text[83] = `CIPHERTEXT_WIDTH'd2741716;
cipher_text[84] = `CIPHERTEXT_WIDTH'd9987937;
cipher_text[85] = `CIPHERTEXT_WIDTH'd13673413;
cipher_text[86] = `CIPHERTEXT_WIDTH'd8392691;
cipher_text[87] = `CIPHERTEXT_WIDTH'd626788;
cipher_text[88] = `CIPHERTEXT_WIDTH'd15916126;
cipher_text[89] = `CIPHERTEXT_WIDTH'd9079298;
cipher_text[90] = `CIPHERTEXT_WIDTH'd5536834;
cipher_text[91] = `CIPHERTEXT_WIDTH'd12076764;
cipher_text[92] = `CIPHERTEXT_WIDTH'd5258654;
cipher_text[93] = `CIPHERTEXT_WIDTH'd13522227;
cipher_text[94] = `CIPHERTEXT_WIDTH'd16627298;
cipher_text[95] = `CIPHERTEXT_WIDTH'd2736894;
cipher_text[96] = `CIPHERTEXT_WIDTH'd8277030;
cipher_text[97] = `CIPHERTEXT_WIDTH'd2805580;
cipher_text[98] = `CIPHERTEXT_WIDTH'd8123467;
cipher_text[99] = `CIPHERTEXT_WIDTH'd5755496;
cipher_text[100] = `CIPHERTEXT_WIDTH'd7593682;
cipher_text[101] = `CIPHERTEXT_WIDTH'd10837940;
cipher_text[102] = `CIPHERTEXT_WIDTH'd13746181;
cipher_text[103] = `CIPHERTEXT_WIDTH'd9394746;
cipher_text[104] = `CIPHERTEXT_WIDTH'd11909383;
cipher_text[105] = `CIPHERTEXT_WIDTH'd13446913;
cipher_text[106] = `CIPHERTEXT_WIDTH'd30769;
cipher_text[107] = `CIPHERTEXT_WIDTH'd15228340;
cipher_text[108] = `CIPHERTEXT_WIDTH'd15843833;
cipher_text[109] = `CIPHERTEXT_WIDTH'd3632983;
cipher_text[110] = `CIPHERTEXT_WIDTH'd4990281;
cipher_text[111] = `CIPHERTEXT_WIDTH'd12563532;
cipher_text[112] = `CIPHERTEXT_WIDTH'd13590773;
cipher_text[113] = `CIPHERTEXT_WIDTH'd2934445;
cipher_text[114] = `CIPHERTEXT_WIDTH'd6601597;
cipher_text[115] = `CIPHERTEXT_WIDTH'd7589383;
cipher_text[116] = `CIPHERTEXT_WIDTH'd7585241;
cipher_text[117] = `CIPHERTEXT_WIDTH'd7277734;
cipher_text[118] = `CIPHERTEXT_WIDTH'd15265425;
cipher_text[119] = `CIPHERTEXT_WIDTH'd13399102;
cipher_text[120] = `CIPHERTEXT_WIDTH'd5914411;
cipher_text[121] = `CIPHERTEXT_WIDTH'd6754255;
cipher_text[122] = `CIPHERTEXT_WIDTH'd15899488;
cipher_text[123] = `CIPHERTEXT_WIDTH'd3389969;
cipher_text[124] = `CIPHERTEXT_WIDTH'd1668206;
cipher_text[125] = `CIPHERTEXT_WIDTH'd15180991;
cipher_text[126] = `CIPHERTEXT_WIDTH'd160085;
cipher_text[127] = `CIPHERTEXT_WIDTH'd5649113;
cipher_text[128] = `CIPHERTEXT_WIDTH'd3826306;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 21;
cipher_text[0] = `CIPHERTEXT_WIDTH'd15646591;
cipher_text[1] = `CIPHERTEXT_WIDTH'd10738127;
cipher_text[2] = `CIPHERTEXT_WIDTH'd214050;
cipher_text[3] = `CIPHERTEXT_WIDTH'd13069250;
cipher_text[4] = `CIPHERTEXT_WIDTH'd12545319;
cipher_text[5] = `CIPHERTEXT_WIDTH'd11323994;
cipher_text[6] = `CIPHERTEXT_WIDTH'd6877121;
cipher_text[7] = `CIPHERTEXT_WIDTH'd1521922;
cipher_text[8] = `CIPHERTEXT_WIDTH'd3986394;
cipher_text[9] = `CIPHERTEXT_WIDTH'd15274289;
cipher_text[10] = `CIPHERTEXT_WIDTH'd15905495;
cipher_text[11] = `CIPHERTEXT_WIDTH'd16058318;
cipher_text[12] = `CIPHERTEXT_WIDTH'd5925219;
cipher_text[13] = `CIPHERTEXT_WIDTH'd12640528;
cipher_text[14] = `CIPHERTEXT_WIDTH'd13515797;
cipher_text[15] = `CIPHERTEXT_WIDTH'd14804200;
cipher_text[16] = `CIPHERTEXT_WIDTH'd4510803;
cipher_text[17] = `CIPHERTEXT_WIDTH'd15461130;
cipher_text[18] = `CIPHERTEXT_WIDTH'd11104078;
cipher_text[19] = `CIPHERTEXT_WIDTH'd15986040;
cipher_text[20] = `CIPHERTEXT_WIDTH'd4890581;
cipher_text[21] = `CIPHERTEXT_WIDTH'd5888795;
cipher_text[22] = `CIPHERTEXT_WIDTH'd4372376;
cipher_text[23] = `CIPHERTEXT_WIDTH'd1606109;
cipher_text[24] = `CIPHERTEXT_WIDTH'd13868714;
cipher_text[25] = `CIPHERTEXT_WIDTH'd3823920;
cipher_text[26] = `CIPHERTEXT_WIDTH'd2246523;
cipher_text[27] = `CIPHERTEXT_WIDTH'd8559192;
cipher_text[28] = `CIPHERTEXT_WIDTH'd6367110;
cipher_text[29] = `CIPHERTEXT_WIDTH'd14627034;
cipher_text[30] = `CIPHERTEXT_WIDTH'd12265398;
cipher_text[31] = `CIPHERTEXT_WIDTH'd6580722;
cipher_text[32] = `CIPHERTEXT_WIDTH'd15791651;
cipher_text[33] = `CIPHERTEXT_WIDTH'd14521098;
cipher_text[34] = `CIPHERTEXT_WIDTH'd14623026;
cipher_text[35] = `CIPHERTEXT_WIDTH'd3957369;
cipher_text[36] = `CIPHERTEXT_WIDTH'd3856744;
cipher_text[37] = `CIPHERTEXT_WIDTH'd7062554;
cipher_text[38] = `CIPHERTEXT_WIDTH'd4941789;
cipher_text[39] = `CIPHERTEXT_WIDTH'd10827642;
cipher_text[40] = `CIPHERTEXT_WIDTH'd3801967;
cipher_text[41] = `CIPHERTEXT_WIDTH'd2274028;
cipher_text[42] = `CIPHERTEXT_WIDTH'd647596;
cipher_text[43] = `CIPHERTEXT_WIDTH'd2602514;
cipher_text[44] = `CIPHERTEXT_WIDTH'd3231606;
cipher_text[45] = `CIPHERTEXT_WIDTH'd14353166;
cipher_text[46] = `CIPHERTEXT_WIDTH'd3971350;
cipher_text[47] = `CIPHERTEXT_WIDTH'd11968411;
cipher_text[48] = `CIPHERTEXT_WIDTH'd4161143;
cipher_text[49] = `CIPHERTEXT_WIDTH'd15252044;
cipher_text[50] = `CIPHERTEXT_WIDTH'd1317912;
cipher_text[51] = `CIPHERTEXT_WIDTH'd16402645;
cipher_text[52] = `CIPHERTEXT_WIDTH'd11196513;
cipher_text[53] = `CIPHERTEXT_WIDTH'd7244240;
cipher_text[54] = `CIPHERTEXT_WIDTH'd14265743;
cipher_text[55] = `CIPHERTEXT_WIDTH'd2765911;
cipher_text[56] = `CIPHERTEXT_WIDTH'd15183625;
cipher_text[57] = `CIPHERTEXT_WIDTH'd8875692;
cipher_text[58] = `CIPHERTEXT_WIDTH'd4273992;
cipher_text[59] = `CIPHERTEXT_WIDTH'd16497789;
cipher_text[60] = `CIPHERTEXT_WIDTH'd2990741;
cipher_text[61] = `CIPHERTEXT_WIDTH'd16023933;
cipher_text[62] = `CIPHERTEXT_WIDTH'd1023496;
cipher_text[63] = `CIPHERTEXT_WIDTH'd4825974;
cipher_text[64] = `CIPHERTEXT_WIDTH'd1434057;
cipher_text[65] = `CIPHERTEXT_WIDTH'd3651892;
cipher_text[66] = `CIPHERTEXT_WIDTH'd14702152;
cipher_text[67] = `CIPHERTEXT_WIDTH'd5513272;
cipher_text[68] = `CIPHERTEXT_WIDTH'd1467126;
cipher_text[69] = `CIPHERTEXT_WIDTH'd15325173;
cipher_text[70] = `CIPHERTEXT_WIDTH'd8426750;
cipher_text[71] = `CIPHERTEXT_WIDTH'd1053028;
cipher_text[72] = `CIPHERTEXT_WIDTH'd5375501;
cipher_text[73] = `CIPHERTEXT_WIDTH'd2707355;
cipher_text[74] = `CIPHERTEXT_WIDTH'd1407380;
cipher_text[75] = `CIPHERTEXT_WIDTH'd15520112;
cipher_text[76] = `CIPHERTEXT_WIDTH'd2779901;
cipher_text[77] = `CIPHERTEXT_WIDTH'd5602005;
cipher_text[78] = `CIPHERTEXT_WIDTH'd16503201;
cipher_text[79] = `CIPHERTEXT_WIDTH'd12299967;
cipher_text[80] = `CIPHERTEXT_WIDTH'd901296;
cipher_text[81] = `CIPHERTEXT_WIDTH'd14112203;
cipher_text[82] = `CIPHERTEXT_WIDTH'd4329743;
cipher_text[83] = `CIPHERTEXT_WIDTH'd7488738;
cipher_text[84] = `CIPHERTEXT_WIDTH'd6644377;
cipher_text[85] = `CIPHERTEXT_WIDTH'd2763295;
cipher_text[86] = `CIPHERTEXT_WIDTH'd8592387;
cipher_text[87] = `CIPHERTEXT_WIDTH'd13148457;
cipher_text[88] = `CIPHERTEXT_WIDTH'd8007259;
cipher_text[89] = `CIPHERTEXT_WIDTH'd7778636;
cipher_text[90] = `CIPHERTEXT_WIDTH'd13237412;
cipher_text[91] = `CIPHERTEXT_WIDTH'd1562316;
cipher_text[92] = `CIPHERTEXT_WIDTH'd9539737;
cipher_text[93] = `CIPHERTEXT_WIDTH'd11416027;
cipher_text[94] = `CIPHERTEXT_WIDTH'd8833831;
cipher_text[95] = `CIPHERTEXT_WIDTH'd13354588;
cipher_text[96] = `CIPHERTEXT_WIDTH'd10273574;
cipher_text[97] = `CIPHERTEXT_WIDTH'd3523271;
cipher_text[98] = `CIPHERTEXT_WIDTH'd11067420;
cipher_text[99] = `CIPHERTEXT_WIDTH'd7249041;
cipher_text[100] = `CIPHERTEXT_WIDTH'd11024473;
cipher_text[101] = `CIPHERTEXT_WIDTH'd12758029;
cipher_text[102] = `CIPHERTEXT_WIDTH'd13294130;
cipher_text[103] = `CIPHERTEXT_WIDTH'd15005380;
cipher_text[104] = `CIPHERTEXT_WIDTH'd3103790;
cipher_text[105] = `CIPHERTEXT_WIDTH'd609749;
cipher_text[106] = `CIPHERTEXT_WIDTH'd7170483;
cipher_text[107] = `CIPHERTEXT_WIDTH'd6520134;
cipher_text[108] = `CIPHERTEXT_WIDTH'd448672;
cipher_text[109] = `CIPHERTEXT_WIDTH'd7520736;
cipher_text[110] = `CIPHERTEXT_WIDTH'd11083117;
cipher_text[111] = `CIPHERTEXT_WIDTH'd2694511;
cipher_text[112] = `CIPHERTEXT_WIDTH'd7094242;
cipher_text[113] = `CIPHERTEXT_WIDTH'd12724434;
cipher_text[114] = `CIPHERTEXT_WIDTH'd8720104;
cipher_text[115] = `CIPHERTEXT_WIDTH'd13865455;
cipher_text[116] = `CIPHERTEXT_WIDTH'd396407;
cipher_text[117] = `CIPHERTEXT_WIDTH'd15577788;
cipher_text[118] = `CIPHERTEXT_WIDTH'd12109798;
cipher_text[119] = `CIPHERTEXT_WIDTH'd9174326;
cipher_text[120] = `CIPHERTEXT_WIDTH'd1794364;
cipher_text[121] = `CIPHERTEXT_WIDTH'd998700;
cipher_text[122] = `CIPHERTEXT_WIDTH'd1620181;
cipher_text[123] = `CIPHERTEXT_WIDTH'd4416866;
cipher_text[124] = `CIPHERTEXT_WIDTH'd9023988;
cipher_text[125] = `CIPHERTEXT_WIDTH'd2254007;
cipher_text[126] = `CIPHERTEXT_WIDTH'd4076205;
cipher_text[127] = `CIPHERTEXT_WIDTH'd1280729;
cipher_text[128] = `CIPHERTEXT_WIDTH'd347006;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 22;
cipher_text[0] = `CIPHERTEXT_WIDTH'd12524981;
cipher_text[1] = `CIPHERTEXT_WIDTH'd4106315;
cipher_text[2] = `CIPHERTEXT_WIDTH'd13074626;
cipher_text[3] = `CIPHERTEXT_WIDTH'd12103190;
cipher_text[4] = `CIPHERTEXT_WIDTH'd7487255;
cipher_text[5] = `CIPHERTEXT_WIDTH'd8405709;
cipher_text[6] = `CIPHERTEXT_WIDTH'd14541616;
cipher_text[7] = `CIPHERTEXT_WIDTH'd603161;
cipher_text[8] = `CIPHERTEXT_WIDTH'd5936108;
cipher_text[9] = `CIPHERTEXT_WIDTH'd3512924;
cipher_text[10] = `CIPHERTEXT_WIDTH'd5718469;
cipher_text[11] = `CIPHERTEXT_WIDTH'd10411243;
cipher_text[12] = `CIPHERTEXT_WIDTH'd1861376;
cipher_text[13] = `CIPHERTEXT_WIDTH'd1124083;
cipher_text[14] = `CIPHERTEXT_WIDTH'd8700183;
cipher_text[15] = `CIPHERTEXT_WIDTH'd16404491;
cipher_text[16] = `CIPHERTEXT_WIDTH'd5283723;
cipher_text[17] = `CIPHERTEXT_WIDTH'd9342540;
cipher_text[18] = `CIPHERTEXT_WIDTH'd15496991;
cipher_text[19] = `CIPHERTEXT_WIDTH'd7102902;
cipher_text[20] = `CIPHERTEXT_WIDTH'd1800719;
cipher_text[21] = `CIPHERTEXT_WIDTH'd7532654;
cipher_text[22] = `CIPHERTEXT_WIDTH'd16226498;
cipher_text[23] = `CIPHERTEXT_WIDTH'd6487610;
cipher_text[24] = `CIPHERTEXT_WIDTH'd599241;
cipher_text[25] = `CIPHERTEXT_WIDTH'd2968265;
cipher_text[26] = `CIPHERTEXT_WIDTH'd8950717;
cipher_text[27] = `CIPHERTEXT_WIDTH'd5642128;
cipher_text[28] = `CIPHERTEXT_WIDTH'd11033679;
cipher_text[29] = `CIPHERTEXT_WIDTH'd7176046;
cipher_text[30] = `CIPHERTEXT_WIDTH'd1802056;
cipher_text[31] = `CIPHERTEXT_WIDTH'd9056478;
cipher_text[32] = `CIPHERTEXT_WIDTH'd9568137;
cipher_text[33] = `CIPHERTEXT_WIDTH'd9082753;
cipher_text[34] = `CIPHERTEXT_WIDTH'd3548554;
cipher_text[35] = `CIPHERTEXT_WIDTH'd7801572;
cipher_text[36] = `CIPHERTEXT_WIDTH'd15349888;
cipher_text[37] = `CIPHERTEXT_WIDTH'd10832114;
cipher_text[38] = `CIPHERTEXT_WIDTH'd9540945;
cipher_text[39] = `CIPHERTEXT_WIDTH'd11826083;
cipher_text[40] = `CIPHERTEXT_WIDTH'd3267292;
cipher_text[41] = `CIPHERTEXT_WIDTH'd12274919;
cipher_text[42] = `CIPHERTEXT_WIDTH'd16140486;
cipher_text[43] = `CIPHERTEXT_WIDTH'd16121196;
cipher_text[44] = `CIPHERTEXT_WIDTH'd1175839;
cipher_text[45] = `CIPHERTEXT_WIDTH'd4954672;
cipher_text[46] = `CIPHERTEXT_WIDTH'd12841034;
cipher_text[47] = `CIPHERTEXT_WIDTH'd6000552;
cipher_text[48] = `CIPHERTEXT_WIDTH'd13507086;
cipher_text[49] = `CIPHERTEXT_WIDTH'd9993504;
cipher_text[50] = `CIPHERTEXT_WIDTH'd9845301;
cipher_text[51] = `CIPHERTEXT_WIDTH'd9702652;
cipher_text[52] = `CIPHERTEXT_WIDTH'd14217393;
cipher_text[53] = `CIPHERTEXT_WIDTH'd3564286;
cipher_text[54] = `CIPHERTEXT_WIDTH'd2888755;
cipher_text[55] = `CIPHERTEXT_WIDTH'd5144061;
cipher_text[56] = `CIPHERTEXT_WIDTH'd10157347;
cipher_text[57] = `CIPHERTEXT_WIDTH'd10697371;
cipher_text[58] = `CIPHERTEXT_WIDTH'd8104880;
cipher_text[59] = `CIPHERTEXT_WIDTH'd6362540;
cipher_text[60] = `CIPHERTEXT_WIDTH'd15028538;
cipher_text[61] = `CIPHERTEXT_WIDTH'd2529378;
cipher_text[62] = `CIPHERTEXT_WIDTH'd15290507;
cipher_text[63] = `CIPHERTEXT_WIDTH'd437418;
cipher_text[64] = `CIPHERTEXT_WIDTH'd7695415;
cipher_text[65] = `CIPHERTEXT_WIDTH'd9099804;
cipher_text[66] = `CIPHERTEXT_WIDTH'd1463412;
cipher_text[67] = `CIPHERTEXT_WIDTH'd15379482;
cipher_text[68] = `CIPHERTEXT_WIDTH'd4034027;
cipher_text[69] = `CIPHERTEXT_WIDTH'd14519790;
cipher_text[70] = `CIPHERTEXT_WIDTH'd13173160;
cipher_text[71] = `CIPHERTEXT_WIDTH'd10808003;
cipher_text[72] = `CIPHERTEXT_WIDTH'd3975305;
cipher_text[73] = `CIPHERTEXT_WIDTH'd11309359;
cipher_text[74] = `CIPHERTEXT_WIDTH'd13278604;
cipher_text[75] = `CIPHERTEXT_WIDTH'd6748102;
cipher_text[76] = `CIPHERTEXT_WIDTH'd3510442;
cipher_text[77] = `CIPHERTEXT_WIDTH'd4170582;
cipher_text[78] = `CIPHERTEXT_WIDTH'd5320062;
cipher_text[79] = `CIPHERTEXT_WIDTH'd10641662;
cipher_text[80] = `CIPHERTEXT_WIDTH'd9196192;
cipher_text[81] = `CIPHERTEXT_WIDTH'd2008272;
cipher_text[82] = `CIPHERTEXT_WIDTH'd14901144;
cipher_text[83] = `CIPHERTEXT_WIDTH'd12643192;
cipher_text[84] = `CIPHERTEXT_WIDTH'd10257054;
cipher_text[85] = `CIPHERTEXT_WIDTH'd6919931;
cipher_text[86] = `CIPHERTEXT_WIDTH'd14144777;
cipher_text[87] = `CIPHERTEXT_WIDTH'd8022869;
cipher_text[88] = `CIPHERTEXT_WIDTH'd5432059;
cipher_text[89] = `CIPHERTEXT_WIDTH'd6922492;
cipher_text[90] = `CIPHERTEXT_WIDTH'd7143346;
cipher_text[91] = `CIPHERTEXT_WIDTH'd531868;
cipher_text[92] = `CIPHERTEXT_WIDTH'd10705703;
cipher_text[93] = `CIPHERTEXT_WIDTH'd13162209;
cipher_text[94] = `CIPHERTEXT_WIDTH'd9654536;
cipher_text[95] = `CIPHERTEXT_WIDTH'd2076496;
cipher_text[96] = `CIPHERTEXT_WIDTH'd14440480;
cipher_text[97] = `CIPHERTEXT_WIDTH'd6515549;
cipher_text[98] = `CIPHERTEXT_WIDTH'd9524166;
cipher_text[99] = `CIPHERTEXT_WIDTH'd3619557;
cipher_text[100] = `CIPHERTEXT_WIDTH'd15481436;
cipher_text[101] = `CIPHERTEXT_WIDTH'd11262080;
cipher_text[102] = `CIPHERTEXT_WIDTH'd6332731;
cipher_text[103] = `CIPHERTEXT_WIDTH'd11399662;
cipher_text[104] = `CIPHERTEXT_WIDTH'd6524622;
cipher_text[105] = `CIPHERTEXT_WIDTH'd3320087;
cipher_text[106] = `CIPHERTEXT_WIDTH'd349555;
cipher_text[107] = `CIPHERTEXT_WIDTH'd13466237;
cipher_text[108] = `CIPHERTEXT_WIDTH'd6451329;
cipher_text[109] = `CIPHERTEXT_WIDTH'd9856175;
cipher_text[110] = `CIPHERTEXT_WIDTH'd14198200;
cipher_text[111] = `CIPHERTEXT_WIDTH'd8215864;
cipher_text[112] = `CIPHERTEXT_WIDTH'd4595606;
cipher_text[113] = `CIPHERTEXT_WIDTH'd301525;
cipher_text[114] = `CIPHERTEXT_WIDTH'd4131143;
cipher_text[115] = `CIPHERTEXT_WIDTH'd15024060;
cipher_text[116] = `CIPHERTEXT_WIDTH'd8572446;
cipher_text[117] = `CIPHERTEXT_WIDTH'd9711552;
cipher_text[118] = `CIPHERTEXT_WIDTH'd15024545;
cipher_text[119] = `CIPHERTEXT_WIDTH'd8680581;
cipher_text[120] = `CIPHERTEXT_WIDTH'd13119792;
cipher_text[121] = `CIPHERTEXT_WIDTH'd12881377;
cipher_text[122] = `CIPHERTEXT_WIDTH'd7740226;
cipher_text[123] = `CIPHERTEXT_WIDTH'd16608245;
cipher_text[124] = `CIPHERTEXT_WIDTH'd6530351;
cipher_text[125] = `CIPHERTEXT_WIDTH'd4177499;
cipher_text[126] = `CIPHERTEXT_WIDTH'd14109197;
cipher_text[127] = `CIPHERTEXT_WIDTH'd5934639;
cipher_text[128] = `CIPHERTEXT_WIDTH'd3550846;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 23;
cipher_text[0] = `CIPHERTEXT_WIDTH'd6664309;
cipher_text[1] = `CIPHERTEXT_WIDTH'd5984974;
cipher_text[2] = `CIPHERTEXT_WIDTH'd1257150;
cipher_text[3] = `CIPHERTEXT_WIDTH'd13965225;
cipher_text[4] = `CIPHERTEXT_WIDTH'd11891398;
cipher_text[5] = `CIPHERTEXT_WIDTH'd4485376;
cipher_text[6] = `CIPHERTEXT_WIDTH'd15057714;
cipher_text[7] = `CIPHERTEXT_WIDTH'd11359997;
cipher_text[8] = `CIPHERTEXT_WIDTH'd15713107;
cipher_text[9] = `CIPHERTEXT_WIDTH'd3502139;
cipher_text[10] = `CIPHERTEXT_WIDTH'd10380442;
cipher_text[11] = `CIPHERTEXT_WIDTH'd1812666;
cipher_text[12] = `CIPHERTEXT_WIDTH'd15870227;
cipher_text[13] = `CIPHERTEXT_WIDTH'd12372227;
cipher_text[14] = `CIPHERTEXT_WIDTH'd2761529;
cipher_text[15] = `CIPHERTEXT_WIDTH'd9063623;
cipher_text[16] = `CIPHERTEXT_WIDTH'd1099834;
cipher_text[17] = `CIPHERTEXT_WIDTH'd5302119;
cipher_text[18] = `CIPHERTEXT_WIDTH'd12018167;
cipher_text[19] = `CIPHERTEXT_WIDTH'd6421825;
cipher_text[20] = `CIPHERTEXT_WIDTH'd1403729;
cipher_text[21] = `CIPHERTEXT_WIDTH'd4686989;
cipher_text[22] = `CIPHERTEXT_WIDTH'd16358737;
cipher_text[23] = `CIPHERTEXT_WIDTH'd15569076;
cipher_text[24] = `CIPHERTEXT_WIDTH'd63834;
cipher_text[25] = `CIPHERTEXT_WIDTH'd3059543;
cipher_text[26] = `CIPHERTEXT_WIDTH'd13665514;
cipher_text[27] = `CIPHERTEXT_WIDTH'd3109156;
cipher_text[28] = `CIPHERTEXT_WIDTH'd14655306;
cipher_text[29] = `CIPHERTEXT_WIDTH'd14209348;
cipher_text[30] = `CIPHERTEXT_WIDTH'd14862387;
cipher_text[31] = `CIPHERTEXT_WIDTH'd14843751;
cipher_text[32] = `CIPHERTEXT_WIDTH'd11735604;
cipher_text[33] = `CIPHERTEXT_WIDTH'd5253610;
cipher_text[34] = `CIPHERTEXT_WIDTH'd16004568;
cipher_text[35] = `CIPHERTEXT_WIDTH'd4257223;
cipher_text[36] = `CIPHERTEXT_WIDTH'd8658079;
cipher_text[37] = `CIPHERTEXT_WIDTH'd4293672;
cipher_text[38] = `CIPHERTEXT_WIDTH'd8073138;
cipher_text[39] = `CIPHERTEXT_WIDTH'd3405779;
cipher_text[40] = `CIPHERTEXT_WIDTH'd1660623;
cipher_text[41] = `CIPHERTEXT_WIDTH'd204996;
cipher_text[42] = `CIPHERTEXT_WIDTH'd6547819;
cipher_text[43] = `CIPHERTEXT_WIDTH'd16130457;
cipher_text[44] = `CIPHERTEXT_WIDTH'd11709204;
cipher_text[45] = `CIPHERTEXT_WIDTH'd12343776;
cipher_text[46] = `CIPHERTEXT_WIDTH'd6488046;
cipher_text[47] = `CIPHERTEXT_WIDTH'd8220318;
cipher_text[48] = `CIPHERTEXT_WIDTH'd10347855;
cipher_text[49] = `CIPHERTEXT_WIDTH'd8430702;
cipher_text[50] = `CIPHERTEXT_WIDTH'd12142747;
cipher_text[51] = `CIPHERTEXT_WIDTH'd8783975;
cipher_text[52] = `CIPHERTEXT_WIDTH'd1608311;
cipher_text[53] = `CIPHERTEXT_WIDTH'd14610575;
cipher_text[54] = `CIPHERTEXT_WIDTH'd14957305;
cipher_text[55] = `CIPHERTEXT_WIDTH'd4365232;
cipher_text[56] = `CIPHERTEXT_WIDTH'd1666932;
cipher_text[57] = `CIPHERTEXT_WIDTH'd11473850;
cipher_text[58] = `CIPHERTEXT_WIDTH'd11643143;
cipher_text[59] = `CIPHERTEXT_WIDTH'd1531605;
cipher_text[60] = `CIPHERTEXT_WIDTH'd7470498;
cipher_text[61] = `CIPHERTEXT_WIDTH'd1315421;
cipher_text[62] = `CIPHERTEXT_WIDTH'd6927387;
cipher_text[63] = `CIPHERTEXT_WIDTH'd7645490;
cipher_text[64] = `CIPHERTEXT_WIDTH'd9857709;
cipher_text[65] = `CIPHERTEXT_WIDTH'd9202818;
cipher_text[66] = `CIPHERTEXT_WIDTH'd12785742;
cipher_text[67] = `CIPHERTEXT_WIDTH'd2463865;
cipher_text[68] = `CIPHERTEXT_WIDTH'd9154758;
cipher_text[69] = `CIPHERTEXT_WIDTH'd11478996;
cipher_text[70] = `CIPHERTEXT_WIDTH'd15984941;
cipher_text[71] = `CIPHERTEXT_WIDTH'd7859436;
cipher_text[72] = `CIPHERTEXT_WIDTH'd4143911;
cipher_text[73] = `CIPHERTEXT_WIDTH'd3990447;
cipher_text[74] = `CIPHERTEXT_WIDTH'd12465139;
cipher_text[75] = `CIPHERTEXT_WIDTH'd12569418;
cipher_text[76] = `CIPHERTEXT_WIDTH'd13149186;
cipher_text[77] = `CIPHERTEXT_WIDTH'd15061817;
cipher_text[78] = `CIPHERTEXT_WIDTH'd16671970;
cipher_text[79] = `CIPHERTEXT_WIDTH'd270093;
cipher_text[80] = `CIPHERTEXT_WIDTH'd13584816;
cipher_text[81] = `CIPHERTEXT_WIDTH'd6451402;
cipher_text[82] = `CIPHERTEXT_WIDTH'd11341059;
cipher_text[83] = `CIPHERTEXT_WIDTH'd8139769;
cipher_text[84] = `CIPHERTEXT_WIDTH'd1922722;
cipher_text[85] = `CIPHERTEXT_WIDTH'd8065342;
cipher_text[86] = `CIPHERTEXT_WIDTH'd1658942;
cipher_text[87] = `CIPHERTEXT_WIDTH'd4250989;
cipher_text[88] = `CIPHERTEXT_WIDTH'd16282472;
cipher_text[89] = `CIPHERTEXT_WIDTH'd16509274;
cipher_text[90] = `CIPHERTEXT_WIDTH'd868060;
cipher_text[91] = `CIPHERTEXT_WIDTH'd15460136;
cipher_text[92] = `CIPHERTEXT_WIDTH'd10841081;
cipher_text[93] = `CIPHERTEXT_WIDTH'd15879800;
cipher_text[94] = `CIPHERTEXT_WIDTH'd14981660;
cipher_text[95] = `CIPHERTEXT_WIDTH'd15209325;
cipher_text[96] = `CIPHERTEXT_WIDTH'd5943840;
cipher_text[97] = `CIPHERTEXT_WIDTH'd5880966;
cipher_text[98] = `CIPHERTEXT_WIDTH'd8523535;
cipher_text[99] = `CIPHERTEXT_WIDTH'd16553735;
cipher_text[100] = `CIPHERTEXT_WIDTH'd1984325;
cipher_text[101] = `CIPHERTEXT_WIDTH'd16297936;
cipher_text[102] = `CIPHERTEXT_WIDTH'd7732906;
cipher_text[103] = `CIPHERTEXT_WIDTH'd1561698;
cipher_text[104] = `CIPHERTEXT_WIDTH'd706822;
cipher_text[105] = `CIPHERTEXT_WIDTH'd6515068;
cipher_text[106] = `CIPHERTEXT_WIDTH'd7218356;
cipher_text[107] = `CIPHERTEXT_WIDTH'd11986679;
cipher_text[108] = `CIPHERTEXT_WIDTH'd16356841;
cipher_text[109] = `CIPHERTEXT_WIDTH'd16547771;
cipher_text[110] = `CIPHERTEXT_WIDTH'd1607289;
cipher_text[111] = `CIPHERTEXT_WIDTH'd10866435;
cipher_text[112] = `CIPHERTEXT_WIDTH'd2219594;
cipher_text[113] = `CIPHERTEXT_WIDTH'd9840127;
cipher_text[114] = `CIPHERTEXT_WIDTH'd2480497;
cipher_text[115] = `CIPHERTEXT_WIDTH'd10445793;
cipher_text[116] = `CIPHERTEXT_WIDTH'd16591221;
cipher_text[117] = `CIPHERTEXT_WIDTH'd12059876;
cipher_text[118] = `CIPHERTEXT_WIDTH'd13674163;
cipher_text[119] = `CIPHERTEXT_WIDTH'd1507816;
cipher_text[120] = `CIPHERTEXT_WIDTH'd11855697;
cipher_text[121] = `CIPHERTEXT_WIDTH'd11257299;
cipher_text[122] = `CIPHERTEXT_WIDTH'd4748145;
cipher_text[123] = `CIPHERTEXT_WIDTH'd3704044;
cipher_text[124] = `CIPHERTEXT_WIDTH'd1808997;
cipher_text[125] = `CIPHERTEXT_WIDTH'd6982263;
cipher_text[126] = `CIPHERTEXT_WIDTH'd505786;
cipher_text[127] = `CIPHERTEXT_WIDTH'd12118038;
cipher_text[128] = `CIPHERTEXT_WIDTH'd6144931;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 24;
cipher_text[0] = `CIPHERTEXT_WIDTH'd4074029;
cipher_text[1] = `CIPHERTEXT_WIDTH'd1063873;
cipher_text[2] = `CIPHERTEXT_WIDTH'd7413118;
cipher_text[3] = `CIPHERTEXT_WIDTH'd8714061;
cipher_text[4] = `CIPHERTEXT_WIDTH'd11047302;
cipher_text[5] = `CIPHERTEXT_WIDTH'd3237739;
cipher_text[6] = `CIPHERTEXT_WIDTH'd7332464;
cipher_text[7] = `CIPHERTEXT_WIDTH'd5542310;
cipher_text[8] = `CIPHERTEXT_WIDTH'd10277041;
cipher_text[9] = `CIPHERTEXT_WIDTH'd12438493;
cipher_text[10] = `CIPHERTEXT_WIDTH'd7267296;
cipher_text[11] = `CIPHERTEXT_WIDTH'd11484553;
cipher_text[12] = `CIPHERTEXT_WIDTH'd11388847;
cipher_text[13] = `CIPHERTEXT_WIDTH'd7645265;
cipher_text[14] = `CIPHERTEXT_WIDTH'd967818;
cipher_text[15] = `CIPHERTEXT_WIDTH'd1282234;
cipher_text[16] = `CIPHERTEXT_WIDTH'd16059436;
cipher_text[17] = `CIPHERTEXT_WIDTH'd14291717;
cipher_text[18] = `CIPHERTEXT_WIDTH'd8945295;
cipher_text[19] = `CIPHERTEXT_WIDTH'd12761932;
cipher_text[20] = `CIPHERTEXT_WIDTH'd9464145;
cipher_text[21] = `CIPHERTEXT_WIDTH'd8427302;
cipher_text[22] = `CIPHERTEXT_WIDTH'd14889738;
cipher_text[23] = `CIPHERTEXT_WIDTH'd10868402;
cipher_text[24] = `CIPHERTEXT_WIDTH'd7985768;
cipher_text[25] = `CIPHERTEXT_WIDTH'd4885480;
cipher_text[26] = `CIPHERTEXT_WIDTH'd7366087;
cipher_text[27] = `CIPHERTEXT_WIDTH'd2576049;
cipher_text[28] = `CIPHERTEXT_WIDTH'd5968008;
cipher_text[29] = `CIPHERTEXT_WIDTH'd13389317;
cipher_text[30] = `CIPHERTEXT_WIDTH'd7889889;
cipher_text[31] = `CIPHERTEXT_WIDTH'd7033089;
cipher_text[32] = `CIPHERTEXT_WIDTH'd9351249;
cipher_text[33] = `CIPHERTEXT_WIDTH'd13706010;
cipher_text[34] = `CIPHERTEXT_WIDTH'd1037984;
cipher_text[35] = `CIPHERTEXT_WIDTH'd6516889;
cipher_text[36] = `CIPHERTEXT_WIDTH'd14674388;
cipher_text[37] = `CIPHERTEXT_WIDTH'd8991240;
cipher_text[38] = `CIPHERTEXT_WIDTH'd14760850;
cipher_text[39] = `CIPHERTEXT_WIDTH'd6075476;
cipher_text[40] = `CIPHERTEXT_WIDTH'd10870951;
cipher_text[41] = `CIPHERTEXT_WIDTH'd1360440;
cipher_text[42] = `CIPHERTEXT_WIDTH'd10084334;
cipher_text[43] = `CIPHERTEXT_WIDTH'd9527648;
cipher_text[44] = `CIPHERTEXT_WIDTH'd15121993;
cipher_text[45] = `CIPHERTEXT_WIDTH'd15718056;
cipher_text[46] = `CIPHERTEXT_WIDTH'd6230088;
cipher_text[47] = `CIPHERTEXT_WIDTH'd9274517;
cipher_text[48] = `CIPHERTEXT_WIDTH'd15659586;
cipher_text[49] = `CIPHERTEXT_WIDTH'd15881832;
cipher_text[50] = `CIPHERTEXT_WIDTH'd4174648;
cipher_text[51] = `CIPHERTEXT_WIDTH'd10950074;
cipher_text[52] = `CIPHERTEXT_WIDTH'd14687556;
cipher_text[53] = `CIPHERTEXT_WIDTH'd11707250;
cipher_text[54] = `CIPHERTEXT_WIDTH'd13367823;
cipher_text[55] = `CIPHERTEXT_WIDTH'd11254444;
cipher_text[56] = `CIPHERTEXT_WIDTH'd412309;
cipher_text[57] = `CIPHERTEXT_WIDTH'd1541102;
cipher_text[58] = `CIPHERTEXT_WIDTH'd4221867;
cipher_text[59] = `CIPHERTEXT_WIDTH'd594903;
cipher_text[60] = `CIPHERTEXT_WIDTH'd2174761;
cipher_text[61] = `CIPHERTEXT_WIDTH'd12341173;
cipher_text[62] = `CIPHERTEXT_WIDTH'd15503602;
cipher_text[63] = `CIPHERTEXT_WIDTH'd5014937;
cipher_text[64] = `CIPHERTEXT_WIDTH'd1876228;
cipher_text[65] = `CIPHERTEXT_WIDTH'd12160497;
cipher_text[66] = `CIPHERTEXT_WIDTH'd10931114;
cipher_text[67] = `CIPHERTEXT_WIDTH'd7143644;
cipher_text[68] = `CIPHERTEXT_WIDTH'd2194708;
cipher_text[69] = `CIPHERTEXT_WIDTH'd11368007;
cipher_text[70] = `CIPHERTEXT_WIDTH'd1776101;
cipher_text[71] = `CIPHERTEXT_WIDTH'd14252755;
cipher_text[72] = `CIPHERTEXT_WIDTH'd2074804;
cipher_text[73] = `CIPHERTEXT_WIDTH'd1373142;
cipher_text[74] = `CIPHERTEXT_WIDTH'd6816;
cipher_text[75] = `CIPHERTEXT_WIDTH'd2233414;
cipher_text[76] = `CIPHERTEXT_WIDTH'd10712147;
cipher_text[77] = `CIPHERTEXT_WIDTH'd3588245;
cipher_text[78] = `CIPHERTEXT_WIDTH'd11743781;
cipher_text[79] = `CIPHERTEXT_WIDTH'd2223355;
cipher_text[80] = `CIPHERTEXT_WIDTH'd5871049;
cipher_text[81] = `CIPHERTEXT_WIDTH'd12989313;
cipher_text[82] = `CIPHERTEXT_WIDTH'd13014252;
cipher_text[83] = `CIPHERTEXT_WIDTH'd3847210;
cipher_text[84] = `CIPHERTEXT_WIDTH'd11478553;
cipher_text[85] = `CIPHERTEXT_WIDTH'd14151061;
cipher_text[86] = `CIPHERTEXT_WIDTH'd2010546;
cipher_text[87] = `CIPHERTEXT_WIDTH'd13144943;
cipher_text[88] = `CIPHERTEXT_WIDTH'd6655408;
cipher_text[89] = `CIPHERTEXT_WIDTH'd4157920;
cipher_text[90] = `CIPHERTEXT_WIDTH'd4561125;
cipher_text[91] = `CIPHERTEXT_WIDTH'd7097742;
cipher_text[92] = `CIPHERTEXT_WIDTH'd7337756;
cipher_text[93] = `CIPHERTEXT_WIDTH'd6114164;
cipher_text[94] = `CIPHERTEXT_WIDTH'd7139220;
cipher_text[95] = `CIPHERTEXT_WIDTH'd11736977;
cipher_text[96] = `CIPHERTEXT_WIDTH'd14038326;
cipher_text[97] = `CIPHERTEXT_WIDTH'd11324273;
cipher_text[98] = `CIPHERTEXT_WIDTH'd16185520;
cipher_text[99] = `CIPHERTEXT_WIDTH'd11807290;
cipher_text[100] = `CIPHERTEXT_WIDTH'd8911039;
cipher_text[101] = `CIPHERTEXT_WIDTH'd2161346;
cipher_text[102] = `CIPHERTEXT_WIDTH'd2080772;
cipher_text[103] = `CIPHERTEXT_WIDTH'd2993897;
cipher_text[104] = `CIPHERTEXT_WIDTH'd13502045;
cipher_text[105] = `CIPHERTEXT_WIDTH'd2791643;
cipher_text[106] = `CIPHERTEXT_WIDTH'd15231211;
cipher_text[107] = `CIPHERTEXT_WIDTH'd2281162;
cipher_text[108] = `CIPHERTEXT_WIDTH'd13018057;
cipher_text[109] = `CIPHERTEXT_WIDTH'd16084582;
cipher_text[110] = `CIPHERTEXT_WIDTH'd10780003;
cipher_text[111] = `CIPHERTEXT_WIDTH'd136248;
cipher_text[112] = `CIPHERTEXT_WIDTH'd1291685;
cipher_text[113] = `CIPHERTEXT_WIDTH'd13409776;
cipher_text[114] = `CIPHERTEXT_WIDTH'd4556542;
cipher_text[115] = `CIPHERTEXT_WIDTH'd16134573;
cipher_text[116] = `CIPHERTEXT_WIDTH'd10915641;
cipher_text[117] = `CIPHERTEXT_WIDTH'd215486;
cipher_text[118] = `CIPHERTEXT_WIDTH'd11815749;
cipher_text[119] = `CIPHERTEXT_WIDTH'd2911231;
cipher_text[120] = `CIPHERTEXT_WIDTH'd7502936;
cipher_text[121] = `CIPHERTEXT_WIDTH'd9022497;
cipher_text[122] = `CIPHERTEXT_WIDTH'd5471953;
cipher_text[123] = `CIPHERTEXT_WIDTH'd16557662;
cipher_text[124] = `CIPHERTEXT_WIDTH'd4793323;
cipher_text[125] = `CIPHERTEXT_WIDTH'd8963511;
cipher_text[126] = `CIPHERTEXT_WIDTH'd4842065;
cipher_text[127] = `CIPHERTEXT_WIDTH'd9078096;
cipher_text[128] = `CIPHERTEXT_WIDTH'd6867393;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 25;
cipher_text[0] = `CIPHERTEXT_WIDTH'd8143962;
cipher_text[1] = `CIPHERTEXT_WIDTH'd14967340;
cipher_text[2] = `CIPHERTEXT_WIDTH'd15876945;
cipher_text[3] = `CIPHERTEXT_WIDTH'd1105745;
cipher_text[4] = `CIPHERTEXT_WIDTH'd2946224;
cipher_text[5] = `CIPHERTEXT_WIDTH'd3177708;
cipher_text[6] = `CIPHERTEXT_WIDTH'd12619054;
cipher_text[7] = `CIPHERTEXT_WIDTH'd8537621;
cipher_text[8] = `CIPHERTEXT_WIDTH'd3397424;
cipher_text[9] = `CIPHERTEXT_WIDTH'd1924917;
cipher_text[10] = `CIPHERTEXT_WIDTH'd15134629;
cipher_text[11] = `CIPHERTEXT_WIDTH'd13837032;
cipher_text[12] = `CIPHERTEXT_WIDTH'd67957;
cipher_text[13] = `CIPHERTEXT_WIDTH'd698718;
cipher_text[14] = `CIPHERTEXT_WIDTH'd9906035;
cipher_text[15] = `CIPHERTEXT_WIDTH'd590481;
cipher_text[16] = `CIPHERTEXT_WIDTH'd5650292;
cipher_text[17] = `CIPHERTEXT_WIDTH'd3790003;
cipher_text[18] = `CIPHERTEXT_WIDTH'd11061515;
cipher_text[19] = `CIPHERTEXT_WIDTH'd16767950;
cipher_text[20] = `CIPHERTEXT_WIDTH'd3272955;
cipher_text[21] = `CIPHERTEXT_WIDTH'd13785690;
cipher_text[22] = `CIPHERTEXT_WIDTH'd10639818;
cipher_text[23] = `CIPHERTEXT_WIDTH'd1182332;
cipher_text[24] = `CIPHERTEXT_WIDTH'd282690;
cipher_text[25] = `CIPHERTEXT_WIDTH'd12225731;
cipher_text[26] = `CIPHERTEXT_WIDTH'd5689169;
cipher_text[27] = `CIPHERTEXT_WIDTH'd440212;
cipher_text[28] = `CIPHERTEXT_WIDTH'd7101675;
cipher_text[29] = `CIPHERTEXT_WIDTH'd13057040;
cipher_text[30] = `CIPHERTEXT_WIDTH'd1952904;
cipher_text[31] = `CIPHERTEXT_WIDTH'd11483902;
cipher_text[32] = `CIPHERTEXT_WIDTH'd12202871;
cipher_text[33] = `CIPHERTEXT_WIDTH'd11914188;
cipher_text[34] = `CIPHERTEXT_WIDTH'd14040936;
cipher_text[35] = `CIPHERTEXT_WIDTH'd1323048;
cipher_text[36] = `CIPHERTEXT_WIDTH'd9344222;
cipher_text[37] = `CIPHERTEXT_WIDTH'd14312139;
cipher_text[38] = `CIPHERTEXT_WIDTH'd6054355;
cipher_text[39] = `CIPHERTEXT_WIDTH'd12522156;
cipher_text[40] = `CIPHERTEXT_WIDTH'd1581764;
cipher_text[41] = `CIPHERTEXT_WIDTH'd10894253;
cipher_text[42] = `CIPHERTEXT_WIDTH'd1775358;
cipher_text[43] = `CIPHERTEXT_WIDTH'd2787457;
cipher_text[44] = `CIPHERTEXT_WIDTH'd3221029;
cipher_text[45] = `CIPHERTEXT_WIDTH'd1032060;
cipher_text[46] = `CIPHERTEXT_WIDTH'd8666514;
cipher_text[47] = `CIPHERTEXT_WIDTH'd13095328;
cipher_text[48] = `CIPHERTEXT_WIDTH'd4228267;
cipher_text[49] = `CIPHERTEXT_WIDTH'd16062538;
cipher_text[50] = `CIPHERTEXT_WIDTH'd8554388;
cipher_text[51] = `CIPHERTEXT_WIDTH'd4460825;
cipher_text[52] = `CIPHERTEXT_WIDTH'd2520104;
cipher_text[53] = `CIPHERTEXT_WIDTH'd10972290;
cipher_text[54] = `CIPHERTEXT_WIDTH'd4230740;
cipher_text[55] = `CIPHERTEXT_WIDTH'd1976548;
cipher_text[56] = `CIPHERTEXT_WIDTH'd16475959;
cipher_text[57] = `CIPHERTEXT_WIDTH'd10722923;
cipher_text[58] = `CIPHERTEXT_WIDTH'd13269474;
cipher_text[59] = `CIPHERTEXT_WIDTH'd10084713;
cipher_text[60] = `CIPHERTEXT_WIDTH'd12001486;
cipher_text[61] = `CIPHERTEXT_WIDTH'd6867069;
cipher_text[62] = `CIPHERTEXT_WIDTH'd12712409;
cipher_text[63] = `CIPHERTEXT_WIDTH'd12294295;
cipher_text[64] = `CIPHERTEXT_WIDTH'd8752002;
cipher_text[65] = `CIPHERTEXT_WIDTH'd14646610;
cipher_text[66] = `CIPHERTEXT_WIDTH'd12079386;
cipher_text[67] = `CIPHERTEXT_WIDTH'd4829726;
cipher_text[68] = `CIPHERTEXT_WIDTH'd13703891;
cipher_text[69] = `CIPHERTEXT_WIDTH'd11361405;
cipher_text[70] = `CIPHERTEXT_WIDTH'd7483845;
cipher_text[71] = `CIPHERTEXT_WIDTH'd8734235;
cipher_text[72] = `CIPHERTEXT_WIDTH'd15246725;
cipher_text[73] = `CIPHERTEXT_WIDTH'd16466145;
cipher_text[74] = `CIPHERTEXT_WIDTH'd9306908;
cipher_text[75] = `CIPHERTEXT_WIDTH'd11544294;
cipher_text[76] = `CIPHERTEXT_WIDTH'd3422488;
cipher_text[77] = `CIPHERTEXT_WIDTH'd6694455;
cipher_text[78] = `CIPHERTEXT_WIDTH'd7183450;
cipher_text[79] = `CIPHERTEXT_WIDTH'd11848241;
cipher_text[80] = `CIPHERTEXT_WIDTH'd12576059;
cipher_text[81] = `CIPHERTEXT_WIDTH'd8778750;
cipher_text[82] = `CIPHERTEXT_WIDTH'd12732762;
cipher_text[83] = `CIPHERTEXT_WIDTH'd12338758;
cipher_text[84] = `CIPHERTEXT_WIDTH'd6481262;
cipher_text[85] = `CIPHERTEXT_WIDTH'd8478580;
cipher_text[86] = `CIPHERTEXT_WIDTH'd8100854;
cipher_text[87] = `CIPHERTEXT_WIDTH'd12629154;
cipher_text[88] = `CIPHERTEXT_WIDTH'd6372711;
cipher_text[89] = `CIPHERTEXT_WIDTH'd10420670;
cipher_text[90] = `CIPHERTEXT_WIDTH'd10310320;
cipher_text[91] = `CIPHERTEXT_WIDTH'd12416035;
cipher_text[92] = `CIPHERTEXT_WIDTH'd382805;
cipher_text[93] = `CIPHERTEXT_WIDTH'd8247290;
cipher_text[94] = `CIPHERTEXT_WIDTH'd8080180;
cipher_text[95] = `CIPHERTEXT_WIDTH'd16157490;
cipher_text[96] = `CIPHERTEXT_WIDTH'd1930228;
cipher_text[97] = `CIPHERTEXT_WIDTH'd15239151;
cipher_text[98] = `CIPHERTEXT_WIDTH'd15723051;
cipher_text[99] = `CIPHERTEXT_WIDTH'd13998539;
cipher_text[100] = `CIPHERTEXT_WIDTH'd16512527;
cipher_text[101] = `CIPHERTEXT_WIDTH'd16588723;
cipher_text[102] = `CIPHERTEXT_WIDTH'd9907560;
cipher_text[103] = `CIPHERTEXT_WIDTH'd16304607;
cipher_text[104] = `CIPHERTEXT_WIDTH'd6576577;
cipher_text[105] = `CIPHERTEXT_WIDTH'd7875254;
cipher_text[106] = `CIPHERTEXT_WIDTH'd5431789;
cipher_text[107] = `CIPHERTEXT_WIDTH'd7673272;
cipher_text[108] = `CIPHERTEXT_WIDTH'd251061;
cipher_text[109] = `CIPHERTEXT_WIDTH'd644042;
cipher_text[110] = `CIPHERTEXT_WIDTH'd952789;
cipher_text[111] = `CIPHERTEXT_WIDTH'd1817098;
cipher_text[112] = `CIPHERTEXT_WIDTH'd4300836;
cipher_text[113] = `CIPHERTEXT_WIDTH'd15365725;
cipher_text[114] = `CIPHERTEXT_WIDTH'd8464660;
cipher_text[115] = `CIPHERTEXT_WIDTH'd14459471;
cipher_text[116] = `CIPHERTEXT_WIDTH'd11719724;
cipher_text[117] = `CIPHERTEXT_WIDTH'd10690709;
cipher_text[118] = `CIPHERTEXT_WIDTH'd7665383;
cipher_text[119] = `CIPHERTEXT_WIDTH'd6365506;
cipher_text[120] = `CIPHERTEXT_WIDTH'd12485498;
cipher_text[121] = `CIPHERTEXT_WIDTH'd6045304;
cipher_text[122] = `CIPHERTEXT_WIDTH'd6540996;
cipher_text[123] = `CIPHERTEXT_WIDTH'd15428742;
cipher_text[124] = `CIPHERTEXT_WIDTH'd2106604;
cipher_text[125] = `CIPHERTEXT_WIDTH'd7677065;
cipher_text[126] = `CIPHERTEXT_WIDTH'd528440;
cipher_text[127] = `CIPHERTEXT_WIDTH'd14852441;
cipher_text[128] = `CIPHERTEXT_WIDTH'd9602945;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 26;
cipher_text[0] = `CIPHERTEXT_WIDTH'd12523673;
cipher_text[1] = `CIPHERTEXT_WIDTH'd528908;
cipher_text[2] = `CIPHERTEXT_WIDTH'd1637390;
cipher_text[3] = `CIPHERTEXT_WIDTH'd9387147;
cipher_text[4] = `CIPHERTEXT_WIDTH'd4178494;
cipher_text[5] = `CIPHERTEXT_WIDTH'd2996131;
cipher_text[6] = `CIPHERTEXT_WIDTH'd7281958;
cipher_text[7] = `CIPHERTEXT_WIDTH'd3055961;
cipher_text[8] = `CIPHERTEXT_WIDTH'd6172839;
cipher_text[9] = `CIPHERTEXT_WIDTH'd6246922;
cipher_text[10] = `CIPHERTEXT_WIDTH'd2875801;
cipher_text[11] = `CIPHERTEXT_WIDTH'd13571372;
cipher_text[12] = `CIPHERTEXT_WIDTH'd515100;
cipher_text[13] = `CIPHERTEXT_WIDTH'd10803835;
cipher_text[14] = `CIPHERTEXT_WIDTH'd2919532;
cipher_text[15] = `CIPHERTEXT_WIDTH'd16399395;
cipher_text[16] = `CIPHERTEXT_WIDTH'd858142;
cipher_text[17] = `CIPHERTEXT_WIDTH'd2218484;
cipher_text[18] = `CIPHERTEXT_WIDTH'd6650420;
cipher_text[19] = `CIPHERTEXT_WIDTH'd5442372;
cipher_text[20] = `CIPHERTEXT_WIDTH'd5553317;
cipher_text[21] = `CIPHERTEXT_WIDTH'd8243205;
cipher_text[22] = `CIPHERTEXT_WIDTH'd11456996;
cipher_text[23] = `CIPHERTEXT_WIDTH'd9143181;
cipher_text[24] = `CIPHERTEXT_WIDTH'd16613244;
cipher_text[25] = `CIPHERTEXT_WIDTH'd8140776;
cipher_text[26] = `CIPHERTEXT_WIDTH'd1857734;
cipher_text[27] = `CIPHERTEXT_WIDTH'd437478;
cipher_text[28] = `CIPHERTEXT_WIDTH'd15273605;
cipher_text[29] = `CIPHERTEXT_WIDTH'd12461704;
cipher_text[30] = `CIPHERTEXT_WIDTH'd7194418;
cipher_text[31] = `CIPHERTEXT_WIDTH'd9649674;
cipher_text[32] = `CIPHERTEXT_WIDTH'd12711695;
cipher_text[33] = `CIPHERTEXT_WIDTH'd625342;
cipher_text[34] = `CIPHERTEXT_WIDTH'd10860528;
cipher_text[35] = `CIPHERTEXT_WIDTH'd7765923;
cipher_text[36] = `CIPHERTEXT_WIDTH'd9401121;
cipher_text[37] = `CIPHERTEXT_WIDTH'd14828557;
cipher_text[38] = `CIPHERTEXT_WIDTH'd5568307;
cipher_text[39] = `CIPHERTEXT_WIDTH'd16426248;
cipher_text[40] = `CIPHERTEXT_WIDTH'd6478289;
cipher_text[41] = `CIPHERTEXT_WIDTH'd6876956;
cipher_text[42] = `CIPHERTEXT_WIDTH'd4007831;
cipher_text[43] = `CIPHERTEXT_WIDTH'd5920431;
cipher_text[44] = `CIPHERTEXT_WIDTH'd310566;
cipher_text[45] = `CIPHERTEXT_WIDTH'd10498136;
cipher_text[46] = `CIPHERTEXT_WIDTH'd9119057;
cipher_text[47] = `CIPHERTEXT_WIDTH'd15984003;
cipher_text[48] = `CIPHERTEXT_WIDTH'd11192252;
cipher_text[49] = `CIPHERTEXT_WIDTH'd16245793;
cipher_text[50] = `CIPHERTEXT_WIDTH'd8031273;
cipher_text[51] = `CIPHERTEXT_WIDTH'd14424621;
cipher_text[52] = `CIPHERTEXT_WIDTH'd1717951;
cipher_text[53] = `CIPHERTEXT_WIDTH'd10858358;
cipher_text[54] = `CIPHERTEXT_WIDTH'd2664373;
cipher_text[55] = `CIPHERTEXT_WIDTH'd5385487;
cipher_text[56] = `CIPHERTEXT_WIDTH'd10126940;
cipher_text[57] = `CIPHERTEXT_WIDTH'd8703584;
cipher_text[58] = `CIPHERTEXT_WIDTH'd1198264;
cipher_text[59] = `CIPHERTEXT_WIDTH'd6750676;
cipher_text[60] = `CIPHERTEXT_WIDTH'd6908827;
cipher_text[61] = `CIPHERTEXT_WIDTH'd4239644;
cipher_text[62] = `CIPHERTEXT_WIDTH'd8454232;
cipher_text[63] = `CIPHERTEXT_WIDTH'd1600061;
cipher_text[64] = `CIPHERTEXT_WIDTH'd4206443;
cipher_text[65] = `CIPHERTEXT_WIDTH'd9103277;
cipher_text[66] = `CIPHERTEXT_WIDTH'd2322707;
cipher_text[67] = `CIPHERTEXT_WIDTH'd563399;
cipher_text[68] = `CIPHERTEXT_WIDTH'd8127617;
cipher_text[69] = `CIPHERTEXT_WIDTH'd10055284;
cipher_text[70] = `CIPHERTEXT_WIDTH'd13256420;
cipher_text[71] = `CIPHERTEXT_WIDTH'd15049485;
cipher_text[72] = `CIPHERTEXT_WIDTH'd3768013;
cipher_text[73] = `CIPHERTEXT_WIDTH'd4273668;
cipher_text[74] = `CIPHERTEXT_WIDTH'd12808091;
cipher_text[75] = `CIPHERTEXT_WIDTH'd7745348;
cipher_text[76] = `CIPHERTEXT_WIDTH'd8728055;
cipher_text[77] = `CIPHERTEXT_WIDTH'd10662622;
cipher_text[78] = `CIPHERTEXT_WIDTH'd11798745;
cipher_text[79] = `CIPHERTEXT_WIDTH'd977539;
cipher_text[80] = `CIPHERTEXT_WIDTH'd9427902;
cipher_text[81] = `CIPHERTEXT_WIDTH'd356712;
cipher_text[82] = `CIPHERTEXT_WIDTH'd7324129;
cipher_text[83] = `CIPHERTEXT_WIDTH'd10694979;
cipher_text[84] = `CIPHERTEXT_WIDTH'd6759790;
cipher_text[85] = `CIPHERTEXT_WIDTH'd9108516;
cipher_text[86] = `CIPHERTEXT_WIDTH'd8424259;
cipher_text[87] = `CIPHERTEXT_WIDTH'd15973031;
cipher_text[88] = `CIPHERTEXT_WIDTH'd8896105;
cipher_text[89] = `CIPHERTEXT_WIDTH'd7906551;
cipher_text[90] = `CIPHERTEXT_WIDTH'd793998;
cipher_text[91] = `CIPHERTEXT_WIDTH'd11792611;
cipher_text[92] = `CIPHERTEXT_WIDTH'd5676732;
cipher_text[93] = `CIPHERTEXT_WIDTH'd6205319;
cipher_text[94] = `CIPHERTEXT_WIDTH'd7966182;
cipher_text[95] = `CIPHERTEXT_WIDTH'd7597455;
cipher_text[96] = `CIPHERTEXT_WIDTH'd4160273;
cipher_text[97] = `CIPHERTEXT_WIDTH'd15921384;
cipher_text[98] = `CIPHERTEXT_WIDTH'd6925795;
cipher_text[99] = `CIPHERTEXT_WIDTH'd1027666;
cipher_text[100] = `CIPHERTEXT_WIDTH'd14193008;
cipher_text[101] = `CIPHERTEXT_WIDTH'd1808318;
cipher_text[102] = `CIPHERTEXT_WIDTH'd1654119;
cipher_text[103] = `CIPHERTEXT_WIDTH'd7138394;
cipher_text[104] = `CIPHERTEXT_WIDTH'd15377615;
cipher_text[105] = `CIPHERTEXT_WIDTH'd2159070;
cipher_text[106] = `CIPHERTEXT_WIDTH'd3845230;
cipher_text[107] = `CIPHERTEXT_WIDTH'd16044005;
cipher_text[108] = `CIPHERTEXT_WIDTH'd11853323;
cipher_text[109] = `CIPHERTEXT_WIDTH'd8232110;
cipher_text[110] = `CIPHERTEXT_WIDTH'd7502079;
cipher_text[111] = `CIPHERTEXT_WIDTH'd6134480;
cipher_text[112] = `CIPHERTEXT_WIDTH'd15300948;
cipher_text[113] = `CIPHERTEXT_WIDTH'd7142529;
cipher_text[114] = `CIPHERTEXT_WIDTH'd6306440;
cipher_text[115] = `CIPHERTEXT_WIDTH'd7180847;
cipher_text[116] = `CIPHERTEXT_WIDTH'd9981630;
cipher_text[117] = `CIPHERTEXT_WIDTH'd3874439;
cipher_text[118] = `CIPHERTEXT_WIDTH'd1174601;
cipher_text[119] = `CIPHERTEXT_WIDTH'd11208756;
cipher_text[120] = `CIPHERTEXT_WIDTH'd9927325;
cipher_text[121] = `CIPHERTEXT_WIDTH'd11316713;
cipher_text[122] = `CIPHERTEXT_WIDTH'd13447924;
cipher_text[123] = `CIPHERTEXT_WIDTH'd604859;
cipher_text[124] = `CIPHERTEXT_WIDTH'd2903597;
cipher_text[125] = `CIPHERTEXT_WIDTH'd15239233;
cipher_text[126] = `CIPHERTEXT_WIDTH'd2624489;
cipher_text[127] = `CIPHERTEXT_WIDTH'd10516142;
cipher_text[128] = `CIPHERTEXT_WIDTH'd11638760;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 27;
cipher_text[0] = `CIPHERTEXT_WIDTH'd15235297;
cipher_text[1] = `CIPHERTEXT_WIDTH'd6566395;
cipher_text[2] = `CIPHERTEXT_WIDTH'd8107383;
cipher_text[3] = `CIPHERTEXT_WIDTH'd9763947;
cipher_text[4] = `CIPHERTEXT_WIDTH'd9841025;
cipher_text[5] = `CIPHERTEXT_WIDTH'd4856888;
cipher_text[6] = `CIPHERTEXT_WIDTH'd336246;
cipher_text[7] = `CIPHERTEXT_WIDTH'd7436216;
cipher_text[8] = `CIPHERTEXT_WIDTH'd8836543;
cipher_text[9] = `CIPHERTEXT_WIDTH'd14707529;
cipher_text[10] = `CIPHERTEXT_WIDTH'd10168467;
cipher_text[11] = `CIPHERTEXT_WIDTH'd8425380;
cipher_text[12] = `CIPHERTEXT_WIDTH'd11817317;
cipher_text[13] = `CIPHERTEXT_WIDTH'd6365293;
cipher_text[14] = `CIPHERTEXT_WIDTH'd12961080;
cipher_text[15] = `CIPHERTEXT_WIDTH'd12225230;
cipher_text[16] = `CIPHERTEXT_WIDTH'd3872545;
cipher_text[17] = `CIPHERTEXT_WIDTH'd14114581;
cipher_text[18] = `CIPHERTEXT_WIDTH'd12435606;
cipher_text[19] = `CIPHERTEXT_WIDTH'd9283669;
cipher_text[20] = `CIPHERTEXT_WIDTH'd2141396;
cipher_text[21] = `CIPHERTEXT_WIDTH'd2383172;
cipher_text[22] = `CIPHERTEXT_WIDTH'd7673817;
cipher_text[23] = `CIPHERTEXT_WIDTH'd3870317;
cipher_text[24] = `CIPHERTEXT_WIDTH'd4244159;
cipher_text[25] = `CIPHERTEXT_WIDTH'd4174471;
cipher_text[26] = `CIPHERTEXT_WIDTH'd1557977;
cipher_text[27] = `CIPHERTEXT_WIDTH'd4227596;
cipher_text[28] = `CIPHERTEXT_WIDTH'd16289408;
cipher_text[29] = `CIPHERTEXT_WIDTH'd5453422;
cipher_text[30] = `CIPHERTEXT_WIDTH'd15674453;
cipher_text[31] = `CIPHERTEXT_WIDTH'd15718754;
cipher_text[32] = `CIPHERTEXT_WIDTH'd13548774;
cipher_text[33] = `CIPHERTEXT_WIDTH'd15963537;
cipher_text[34] = `CIPHERTEXT_WIDTH'd12772589;
cipher_text[35] = `CIPHERTEXT_WIDTH'd1552159;
cipher_text[36] = `CIPHERTEXT_WIDTH'd14951574;
cipher_text[37] = `CIPHERTEXT_WIDTH'd14959046;
cipher_text[38] = `CIPHERTEXT_WIDTH'd3198057;
cipher_text[39] = `CIPHERTEXT_WIDTH'd11210910;
cipher_text[40] = `CIPHERTEXT_WIDTH'd7589016;
cipher_text[41] = `CIPHERTEXT_WIDTH'd11663213;
cipher_text[42] = `CIPHERTEXT_WIDTH'd4529273;
cipher_text[43] = `CIPHERTEXT_WIDTH'd9304127;
cipher_text[44] = `CIPHERTEXT_WIDTH'd6234106;
cipher_text[45] = `CIPHERTEXT_WIDTH'd13980244;
cipher_text[46] = `CIPHERTEXT_WIDTH'd2962102;
cipher_text[47] = `CIPHERTEXT_WIDTH'd14153453;
cipher_text[48] = `CIPHERTEXT_WIDTH'd16558641;
cipher_text[49] = `CIPHERTEXT_WIDTH'd13285601;
cipher_text[50] = `CIPHERTEXT_WIDTH'd13950957;
cipher_text[51] = `CIPHERTEXT_WIDTH'd6107731;
cipher_text[52] = `CIPHERTEXT_WIDTH'd8399519;
cipher_text[53] = `CIPHERTEXT_WIDTH'd16381051;
cipher_text[54] = `CIPHERTEXT_WIDTH'd5513506;
cipher_text[55] = `CIPHERTEXT_WIDTH'd4749840;
cipher_text[56] = `CIPHERTEXT_WIDTH'd6651071;
cipher_text[57] = `CIPHERTEXT_WIDTH'd16374323;
cipher_text[58] = `CIPHERTEXT_WIDTH'd1005063;
cipher_text[59] = `CIPHERTEXT_WIDTH'd2453604;
cipher_text[60] = `CIPHERTEXT_WIDTH'd16039479;
cipher_text[61] = `CIPHERTEXT_WIDTH'd6009000;
cipher_text[62] = `CIPHERTEXT_WIDTH'd10545774;
cipher_text[63] = `CIPHERTEXT_WIDTH'd1160110;
cipher_text[64] = `CIPHERTEXT_WIDTH'd13807723;
cipher_text[65] = `CIPHERTEXT_WIDTH'd16346220;
cipher_text[66] = `CIPHERTEXT_WIDTH'd4164158;
cipher_text[67] = `CIPHERTEXT_WIDTH'd3498146;
cipher_text[68] = `CIPHERTEXT_WIDTH'd12247264;
cipher_text[69] = `CIPHERTEXT_WIDTH'd13387305;
cipher_text[70] = `CIPHERTEXT_WIDTH'd12992173;
cipher_text[71] = `CIPHERTEXT_WIDTH'd2039423;
cipher_text[72] = `CIPHERTEXT_WIDTH'd8691381;
cipher_text[73] = `CIPHERTEXT_WIDTH'd528253;
cipher_text[74] = `CIPHERTEXT_WIDTH'd1403435;
cipher_text[75] = `CIPHERTEXT_WIDTH'd274687;
cipher_text[76] = `CIPHERTEXT_WIDTH'd8992;
cipher_text[77] = `CIPHERTEXT_WIDTH'd146106;
cipher_text[78] = `CIPHERTEXT_WIDTH'd13934218;
cipher_text[79] = `CIPHERTEXT_WIDTH'd14140692;
cipher_text[80] = `CIPHERTEXT_WIDTH'd9306458;
cipher_text[81] = `CIPHERTEXT_WIDTH'd8501188;
cipher_text[82] = `CIPHERTEXT_WIDTH'd2206607;
cipher_text[83] = `CIPHERTEXT_WIDTH'd6294784;
cipher_text[84] = `CIPHERTEXT_WIDTH'd10101476;
cipher_text[85] = `CIPHERTEXT_WIDTH'd4085870;
cipher_text[86] = `CIPHERTEXT_WIDTH'd1409116;
cipher_text[87] = `CIPHERTEXT_WIDTH'd1929976;
cipher_text[88] = `CIPHERTEXT_WIDTH'd14851046;
cipher_text[89] = `CIPHERTEXT_WIDTH'd2338743;
cipher_text[90] = `CIPHERTEXT_WIDTH'd14831511;
cipher_text[91] = `CIPHERTEXT_WIDTH'd12168942;
cipher_text[92] = `CIPHERTEXT_WIDTH'd14623431;
cipher_text[93] = `CIPHERTEXT_WIDTH'd5118713;
cipher_text[94] = `CIPHERTEXT_WIDTH'd11599563;
cipher_text[95] = `CIPHERTEXT_WIDTH'd1398289;
cipher_text[96] = `CIPHERTEXT_WIDTH'd15496186;
cipher_text[97] = `CIPHERTEXT_WIDTH'd3930321;
cipher_text[98] = `CIPHERTEXT_WIDTH'd8062096;
cipher_text[99] = `CIPHERTEXT_WIDTH'd5709817;
cipher_text[100] = `CIPHERTEXT_WIDTH'd2359222;
cipher_text[101] = `CIPHERTEXT_WIDTH'd9349381;
cipher_text[102] = `CIPHERTEXT_WIDTH'd148811;
cipher_text[103] = `CIPHERTEXT_WIDTH'd9869675;
cipher_text[104] = `CIPHERTEXT_WIDTH'd429032;
cipher_text[105] = `CIPHERTEXT_WIDTH'd14865033;
cipher_text[106] = `CIPHERTEXT_WIDTH'd3735555;
cipher_text[107] = `CIPHERTEXT_WIDTH'd8078540;
cipher_text[108] = `CIPHERTEXT_WIDTH'd2464290;
cipher_text[109] = `CIPHERTEXT_WIDTH'd2472212;
cipher_text[110] = `CIPHERTEXT_WIDTH'd4491111;
cipher_text[111] = `CIPHERTEXT_WIDTH'd1024374;
cipher_text[112] = `CIPHERTEXT_WIDTH'd2124905;
cipher_text[113] = `CIPHERTEXT_WIDTH'd7921966;
cipher_text[114] = `CIPHERTEXT_WIDTH'd8918607;
cipher_text[115] = `CIPHERTEXT_WIDTH'd10696521;
cipher_text[116] = `CIPHERTEXT_WIDTH'd10857407;
cipher_text[117] = `CIPHERTEXT_WIDTH'd735459;
cipher_text[118] = `CIPHERTEXT_WIDTH'd7348189;
cipher_text[119] = `CIPHERTEXT_WIDTH'd3326268;
cipher_text[120] = `CIPHERTEXT_WIDTH'd11999667;
cipher_text[121] = `CIPHERTEXT_WIDTH'd16084158;
cipher_text[122] = `CIPHERTEXT_WIDTH'd9005615;
cipher_text[123] = `CIPHERTEXT_WIDTH'd14161216;
cipher_text[124] = `CIPHERTEXT_WIDTH'd10831885;
cipher_text[125] = `CIPHERTEXT_WIDTH'd8671097;
cipher_text[126] = `CIPHERTEXT_WIDTH'd627633;
cipher_text[127] = `CIPHERTEXT_WIDTH'd13715934;
cipher_text[128] = `CIPHERTEXT_WIDTH'd9381824;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 28;
cipher_text[0] = `CIPHERTEXT_WIDTH'd164103;
cipher_text[1] = `CIPHERTEXT_WIDTH'd4819319;
cipher_text[2] = `CIPHERTEXT_WIDTH'd11029653;
cipher_text[3] = `CIPHERTEXT_WIDTH'd9749661;
cipher_text[4] = `CIPHERTEXT_WIDTH'd5403844;
cipher_text[5] = `CIPHERTEXT_WIDTH'd7112197;
cipher_text[6] = `CIPHERTEXT_WIDTH'd8091668;
cipher_text[7] = `CIPHERTEXT_WIDTH'd9644763;
cipher_text[8] = `CIPHERTEXT_WIDTH'd8923014;
cipher_text[9] = `CIPHERTEXT_WIDTH'd5130948;
cipher_text[10] = `CIPHERTEXT_WIDTH'd11736715;
cipher_text[11] = `CIPHERTEXT_WIDTH'd576798;
cipher_text[12] = `CIPHERTEXT_WIDTH'd4452128;
cipher_text[13] = `CIPHERTEXT_WIDTH'd3475935;
cipher_text[14] = `CIPHERTEXT_WIDTH'd7213020;
cipher_text[15] = `CIPHERTEXT_WIDTH'd13060132;
cipher_text[16] = `CIPHERTEXT_WIDTH'd10155642;
cipher_text[17] = `CIPHERTEXT_WIDTH'd542766;
cipher_text[18] = `CIPHERTEXT_WIDTH'd5033501;
cipher_text[19] = `CIPHERTEXT_WIDTH'd11028782;
cipher_text[20] = `CIPHERTEXT_WIDTH'd4727392;
cipher_text[21] = `CIPHERTEXT_WIDTH'd16144918;
cipher_text[22] = `CIPHERTEXT_WIDTH'd4112552;
cipher_text[23] = `CIPHERTEXT_WIDTH'd3062197;
cipher_text[24] = `CIPHERTEXT_WIDTH'd3691092;
cipher_text[25] = `CIPHERTEXT_WIDTH'd11644918;
cipher_text[26] = `CIPHERTEXT_WIDTH'd12786582;
cipher_text[27] = `CIPHERTEXT_WIDTH'd6232311;
cipher_text[28] = `CIPHERTEXT_WIDTH'd2852355;
cipher_text[29] = `CIPHERTEXT_WIDTH'd1829516;
cipher_text[30] = `CIPHERTEXT_WIDTH'd8816388;
cipher_text[31] = `CIPHERTEXT_WIDTH'd7683441;
cipher_text[32] = `CIPHERTEXT_WIDTH'd14076980;
cipher_text[33] = `CIPHERTEXT_WIDTH'd15274719;
cipher_text[34] = `CIPHERTEXT_WIDTH'd7848966;
cipher_text[35] = `CIPHERTEXT_WIDTH'd15569812;
cipher_text[36] = `CIPHERTEXT_WIDTH'd8976802;
cipher_text[37] = `CIPHERTEXT_WIDTH'd12517227;
cipher_text[38] = `CIPHERTEXT_WIDTH'd247272;
cipher_text[39] = `CIPHERTEXT_WIDTH'd938243;
cipher_text[40] = `CIPHERTEXT_WIDTH'd10099912;
cipher_text[41] = `CIPHERTEXT_WIDTH'd7374806;
cipher_text[42] = `CIPHERTEXT_WIDTH'd4208079;
cipher_text[43] = `CIPHERTEXT_WIDTH'd355785;
cipher_text[44] = `CIPHERTEXT_WIDTH'd2153201;
cipher_text[45] = `CIPHERTEXT_WIDTH'd13737165;
cipher_text[46] = `CIPHERTEXT_WIDTH'd15218086;
cipher_text[47] = `CIPHERTEXT_WIDTH'd2089021;
cipher_text[48] = `CIPHERTEXT_WIDTH'd3219147;
cipher_text[49] = `CIPHERTEXT_WIDTH'd7953366;
cipher_text[50] = `CIPHERTEXT_WIDTH'd594793;
cipher_text[51] = `CIPHERTEXT_WIDTH'd9960327;
cipher_text[52] = `CIPHERTEXT_WIDTH'd2922496;
cipher_text[53] = `CIPHERTEXT_WIDTH'd5615919;
cipher_text[54] = `CIPHERTEXT_WIDTH'd4201829;
cipher_text[55] = `CIPHERTEXT_WIDTH'd15370466;
cipher_text[56] = `CIPHERTEXT_WIDTH'd13394745;
cipher_text[57] = `CIPHERTEXT_WIDTH'd8965362;
cipher_text[58] = `CIPHERTEXT_WIDTH'd4564383;
cipher_text[59] = `CIPHERTEXT_WIDTH'd13329039;
cipher_text[60] = `CIPHERTEXT_WIDTH'd264579;
cipher_text[61] = `CIPHERTEXT_WIDTH'd4274049;
cipher_text[62] = `CIPHERTEXT_WIDTH'd15132934;
cipher_text[63] = `CIPHERTEXT_WIDTH'd7801658;
cipher_text[64] = `CIPHERTEXT_WIDTH'd11088758;
cipher_text[65] = `CIPHERTEXT_WIDTH'd14248666;
cipher_text[66] = `CIPHERTEXT_WIDTH'd1079113;
cipher_text[67] = `CIPHERTEXT_WIDTH'd7127909;
cipher_text[68] = `CIPHERTEXT_WIDTH'd13341669;
cipher_text[69] = `CIPHERTEXT_WIDTH'd16177161;
cipher_text[70] = `CIPHERTEXT_WIDTH'd10897140;
cipher_text[71] = `CIPHERTEXT_WIDTH'd14108790;
cipher_text[72] = `CIPHERTEXT_WIDTH'd4456800;
cipher_text[73] = `CIPHERTEXT_WIDTH'd10776704;
cipher_text[74] = `CIPHERTEXT_WIDTH'd7832053;
cipher_text[75] = `CIPHERTEXT_WIDTH'd7805546;
cipher_text[76] = `CIPHERTEXT_WIDTH'd16614105;
cipher_text[77] = `CIPHERTEXT_WIDTH'd3444003;
cipher_text[78] = `CIPHERTEXT_WIDTH'd10078429;
cipher_text[79] = `CIPHERTEXT_WIDTH'd8125071;
cipher_text[80] = `CIPHERTEXT_WIDTH'd2700087;
cipher_text[81] = `CIPHERTEXT_WIDTH'd3260403;
cipher_text[82] = `CIPHERTEXT_WIDTH'd11207144;
cipher_text[83] = `CIPHERTEXT_WIDTH'd15121987;
cipher_text[84] = `CIPHERTEXT_WIDTH'd4702664;
cipher_text[85] = `CIPHERTEXT_WIDTH'd9148938;
cipher_text[86] = `CIPHERTEXT_WIDTH'd5070249;
cipher_text[87] = `CIPHERTEXT_WIDTH'd5088378;
cipher_text[88] = `CIPHERTEXT_WIDTH'd12954383;
cipher_text[89] = `CIPHERTEXT_WIDTH'd6622945;
cipher_text[90] = `CIPHERTEXT_WIDTH'd16505661;
cipher_text[91] = `CIPHERTEXT_WIDTH'd6972408;
cipher_text[92] = `CIPHERTEXT_WIDTH'd11105371;
cipher_text[93] = `CIPHERTEXT_WIDTH'd8663293;
cipher_text[94] = `CIPHERTEXT_WIDTH'd1108878;
cipher_text[95] = `CIPHERTEXT_WIDTH'd8257619;
cipher_text[96] = `CIPHERTEXT_WIDTH'd9420314;
cipher_text[97] = `CIPHERTEXT_WIDTH'd6131942;
cipher_text[98] = `CIPHERTEXT_WIDTH'd8679628;
cipher_text[99] = `CIPHERTEXT_WIDTH'd7185344;
cipher_text[100] = `CIPHERTEXT_WIDTH'd2703141;
cipher_text[101] = `CIPHERTEXT_WIDTH'd892889;
cipher_text[102] = `CIPHERTEXT_WIDTH'd13907818;
cipher_text[103] = `CIPHERTEXT_WIDTH'd11770292;
cipher_text[104] = `CIPHERTEXT_WIDTH'd3792024;
cipher_text[105] = `CIPHERTEXT_WIDTH'd12749802;
cipher_text[106] = `CIPHERTEXT_WIDTH'd8224528;
cipher_text[107] = `CIPHERTEXT_WIDTH'd7016875;
cipher_text[108] = `CIPHERTEXT_WIDTH'd14662278;
cipher_text[109] = `CIPHERTEXT_WIDTH'd6919015;
cipher_text[110] = `CIPHERTEXT_WIDTH'd15499267;
cipher_text[111] = `CIPHERTEXT_WIDTH'd12477479;
cipher_text[112] = `CIPHERTEXT_WIDTH'd12201387;
cipher_text[113] = `CIPHERTEXT_WIDTH'd12322564;
cipher_text[114] = `CIPHERTEXT_WIDTH'd4724652;
cipher_text[115] = `CIPHERTEXT_WIDTH'd8946104;
cipher_text[116] = `CIPHERTEXT_WIDTH'd10346812;
cipher_text[117] = `CIPHERTEXT_WIDTH'd6426292;
cipher_text[118] = `CIPHERTEXT_WIDTH'd5577467;
cipher_text[119] = `CIPHERTEXT_WIDTH'd16453390;
cipher_text[120] = `CIPHERTEXT_WIDTH'd7388291;
cipher_text[121] = `CIPHERTEXT_WIDTH'd2393686;
cipher_text[122] = `CIPHERTEXT_WIDTH'd7065496;
cipher_text[123] = `CIPHERTEXT_WIDTH'd13047563;
cipher_text[124] = `CIPHERTEXT_WIDTH'd11845690;
cipher_text[125] = `CIPHERTEXT_WIDTH'd1194754;
cipher_text[126] = `CIPHERTEXT_WIDTH'd7935417;
cipher_text[127] = `CIPHERTEXT_WIDTH'd16697290;
cipher_text[128] = `CIPHERTEXT_WIDTH'd4299461;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 29;
cipher_text[0] = `CIPHERTEXT_WIDTH'd16770478;
cipher_text[1] = `CIPHERTEXT_WIDTH'd2415432;
cipher_text[2] = `CIPHERTEXT_WIDTH'd11986233;
cipher_text[3] = `CIPHERTEXT_WIDTH'd7345977;
cipher_text[4] = `CIPHERTEXT_WIDTH'd2066016;
cipher_text[5] = `CIPHERTEXT_WIDTH'd2827824;
cipher_text[6] = `CIPHERTEXT_WIDTH'd2366060;
cipher_text[7] = `CIPHERTEXT_WIDTH'd808122;
cipher_text[8] = `CIPHERTEXT_WIDTH'd12615322;
cipher_text[9] = `CIPHERTEXT_WIDTH'd7150127;
cipher_text[10] = `CIPHERTEXT_WIDTH'd10640916;
cipher_text[11] = `CIPHERTEXT_WIDTH'd6965270;
cipher_text[12] = `CIPHERTEXT_WIDTH'd2441054;
cipher_text[13] = `CIPHERTEXT_WIDTH'd7715294;
cipher_text[14] = `CIPHERTEXT_WIDTH'd13645915;
cipher_text[15] = `CIPHERTEXT_WIDTH'd9905790;
cipher_text[16] = `CIPHERTEXT_WIDTH'd2138647;
cipher_text[17] = `CIPHERTEXT_WIDTH'd4846151;
cipher_text[18] = `CIPHERTEXT_WIDTH'd14589415;
cipher_text[19] = `CIPHERTEXT_WIDTH'd13990473;
cipher_text[20] = `CIPHERTEXT_WIDTH'd12878423;
cipher_text[21] = `CIPHERTEXT_WIDTH'd6030680;
cipher_text[22] = `CIPHERTEXT_WIDTH'd6415401;
cipher_text[23] = `CIPHERTEXT_WIDTH'd9755424;
cipher_text[24] = `CIPHERTEXT_WIDTH'd5291039;
cipher_text[25] = `CIPHERTEXT_WIDTH'd3833518;
cipher_text[26] = `CIPHERTEXT_WIDTH'd13111187;
cipher_text[27] = `CIPHERTEXT_WIDTH'd15090548;
cipher_text[28] = `CIPHERTEXT_WIDTH'd5227100;
cipher_text[29] = `CIPHERTEXT_WIDTH'd4088571;
cipher_text[30] = `CIPHERTEXT_WIDTH'd12319378;
cipher_text[31] = `CIPHERTEXT_WIDTH'd14625178;
cipher_text[32] = `CIPHERTEXT_WIDTH'd8246783;
cipher_text[33] = `CIPHERTEXT_WIDTH'd4763705;
cipher_text[34] = `CIPHERTEXT_WIDTH'd2635844;
cipher_text[35] = `CIPHERTEXT_WIDTH'd13359647;
cipher_text[36] = `CIPHERTEXT_WIDTH'd12394551;
cipher_text[37] = `CIPHERTEXT_WIDTH'd4301403;
cipher_text[38] = `CIPHERTEXT_WIDTH'd8437581;
cipher_text[39] = `CIPHERTEXT_WIDTH'd4823407;
cipher_text[40] = `CIPHERTEXT_WIDTH'd9435035;
cipher_text[41] = `CIPHERTEXT_WIDTH'd14616107;
cipher_text[42] = `CIPHERTEXT_WIDTH'd6536812;
cipher_text[43] = `CIPHERTEXT_WIDTH'd12658803;
cipher_text[44] = `CIPHERTEXT_WIDTH'd7508572;
cipher_text[45] = `CIPHERTEXT_WIDTH'd16203466;
cipher_text[46] = `CIPHERTEXT_WIDTH'd10749971;
cipher_text[47] = `CIPHERTEXT_WIDTH'd6974084;
cipher_text[48] = `CIPHERTEXT_WIDTH'd16434171;
cipher_text[49] = `CIPHERTEXT_WIDTH'd13483701;
cipher_text[50] = `CIPHERTEXT_WIDTH'd4590045;
cipher_text[51] = `CIPHERTEXT_WIDTH'd14365283;
cipher_text[52] = `CIPHERTEXT_WIDTH'd9932123;
cipher_text[53] = `CIPHERTEXT_WIDTH'd13628459;
cipher_text[54] = `CIPHERTEXT_WIDTH'd14910616;
cipher_text[55] = `CIPHERTEXT_WIDTH'd3808184;
cipher_text[56] = `CIPHERTEXT_WIDTH'd5805878;
cipher_text[57] = `CIPHERTEXT_WIDTH'd12668195;
cipher_text[58] = `CIPHERTEXT_WIDTH'd5462311;
cipher_text[59] = `CIPHERTEXT_WIDTH'd2697919;
cipher_text[60] = `CIPHERTEXT_WIDTH'd15496610;
cipher_text[61] = `CIPHERTEXT_WIDTH'd12994152;
cipher_text[62] = `CIPHERTEXT_WIDTH'd10089073;
cipher_text[63] = `CIPHERTEXT_WIDTH'd12155833;
cipher_text[64] = `CIPHERTEXT_WIDTH'd804189;
cipher_text[65] = `CIPHERTEXT_WIDTH'd16168515;
cipher_text[66] = `CIPHERTEXT_WIDTH'd8791401;
cipher_text[67] = `CIPHERTEXT_WIDTH'd6053626;
cipher_text[68] = `CIPHERTEXT_WIDTH'd9062907;
cipher_text[69] = `CIPHERTEXT_WIDTH'd14999394;
cipher_text[70] = `CIPHERTEXT_WIDTH'd15591866;
cipher_text[71] = `CIPHERTEXT_WIDTH'd7055911;
cipher_text[72] = `CIPHERTEXT_WIDTH'd4677619;
cipher_text[73] = `CIPHERTEXT_WIDTH'd16263268;
cipher_text[74] = `CIPHERTEXT_WIDTH'd8680705;
cipher_text[75] = `CIPHERTEXT_WIDTH'd6785419;
cipher_text[76] = `CIPHERTEXT_WIDTH'd2798883;
cipher_text[77] = `CIPHERTEXT_WIDTH'd14853109;
cipher_text[78] = `CIPHERTEXT_WIDTH'd2930215;
cipher_text[79] = `CIPHERTEXT_WIDTH'd6148855;
cipher_text[80] = `CIPHERTEXT_WIDTH'd2317457;
cipher_text[81] = `CIPHERTEXT_WIDTH'd1180689;
cipher_text[82] = `CIPHERTEXT_WIDTH'd13385209;
cipher_text[83] = `CIPHERTEXT_WIDTH'd11707052;
cipher_text[84] = `CIPHERTEXT_WIDTH'd5005828;
cipher_text[85] = `CIPHERTEXT_WIDTH'd16119056;
cipher_text[86] = `CIPHERTEXT_WIDTH'd1766754;
cipher_text[87] = `CIPHERTEXT_WIDTH'd3892138;
cipher_text[88] = `CIPHERTEXT_WIDTH'd9030123;
cipher_text[89] = `CIPHERTEXT_WIDTH'd8981583;
cipher_text[90] = `CIPHERTEXT_WIDTH'd12808853;
cipher_text[91] = `CIPHERTEXT_WIDTH'd1925150;
cipher_text[92] = `CIPHERTEXT_WIDTH'd13093098;
cipher_text[93] = `CIPHERTEXT_WIDTH'd12471035;
cipher_text[94] = `CIPHERTEXT_WIDTH'd10943561;
cipher_text[95] = `CIPHERTEXT_WIDTH'd8313096;
cipher_text[96] = `CIPHERTEXT_WIDTH'd9362173;
cipher_text[97] = `CIPHERTEXT_WIDTH'd3261917;
cipher_text[98] = `CIPHERTEXT_WIDTH'd9701848;
cipher_text[99] = `CIPHERTEXT_WIDTH'd6673793;
cipher_text[100] = `CIPHERTEXT_WIDTH'd16146148;
cipher_text[101] = `CIPHERTEXT_WIDTH'd10270640;
cipher_text[102] = `CIPHERTEXT_WIDTH'd7512214;
cipher_text[103] = `CIPHERTEXT_WIDTH'd3534718;
cipher_text[104] = `CIPHERTEXT_WIDTH'd3461947;
cipher_text[105] = `CIPHERTEXT_WIDTH'd9618207;
cipher_text[106] = `CIPHERTEXT_WIDTH'd3098841;
cipher_text[107] = `CIPHERTEXT_WIDTH'd3694281;
cipher_text[108] = `CIPHERTEXT_WIDTH'd15446308;
cipher_text[109] = `CIPHERTEXT_WIDTH'd3618827;
cipher_text[110] = `CIPHERTEXT_WIDTH'd15959366;
cipher_text[111] = `CIPHERTEXT_WIDTH'd9804407;
cipher_text[112] = `CIPHERTEXT_WIDTH'd6886981;
cipher_text[113] = `CIPHERTEXT_WIDTH'd14827346;
cipher_text[114] = `CIPHERTEXT_WIDTH'd11278896;
cipher_text[115] = `CIPHERTEXT_WIDTH'd11540450;
cipher_text[116] = `CIPHERTEXT_WIDTH'd16271194;
cipher_text[117] = `CIPHERTEXT_WIDTH'd2738215;
cipher_text[118] = `CIPHERTEXT_WIDTH'd5354192;
cipher_text[119] = `CIPHERTEXT_WIDTH'd13047900;
cipher_text[120] = `CIPHERTEXT_WIDTH'd6064082;
cipher_text[121] = `CIPHERTEXT_WIDTH'd3871778;
cipher_text[122] = `CIPHERTEXT_WIDTH'd8756424;
cipher_text[123] = `CIPHERTEXT_WIDTH'd9403105;
cipher_text[124] = `CIPHERTEXT_WIDTH'd8446140;
cipher_text[125] = `CIPHERTEXT_WIDTH'd5547219;
cipher_text[126] = `CIPHERTEXT_WIDTH'd115330;
cipher_text[127] = `CIPHERTEXT_WIDTH'd15428927;
cipher_text[128] = `CIPHERTEXT_WIDTH'd2575035;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 30;
cipher_text[0] = `CIPHERTEXT_WIDTH'd13955836;
cipher_text[1] = `CIPHERTEXT_WIDTH'd10848619;
cipher_text[2] = `CIPHERTEXT_WIDTH'd6258604;
cipher_text[3] = `CIPHERTEXT_WIDTH'd12870306;
cipher_text[4] = `CIPHERTEXT_WIDTH'd1003477;
cipher_text[5] = `CIPHERTEXT_WIDTH'd9664969;
cipher_text[6] = `CIPHERTEXT_WIDTH'd16248217;
cipher_text[7] = `CIPHERTEXT_WIDTH'd13904564;
cipher_text[8] = `CIPHERTEXT_WIDTH'd1011147;
cipher_text[9] = `CIPHERTEXT_WIDTH'd11581612;
cipher_text[10] = `CIPHERTEXT_WIDTH'd14459610;
cipher_text[11] = `CIPHERTEXT_WIDTH'd4811148;
cipher_text[12] = `CIPHERTEXT_WIDTH'd10382086;
cipher_text[13] = `CIPHERTEXT_WIDTH'd11615023;
cipher_text[14] = `CIPHERTEXT_WIDTH'd4406115;
cipher_text[15] = `CIPHERTEXT_WIDTH'd9535997;
cipher_text[16] = `CIPHERTEXT_WIDTH'd14383081;
cipher_text[17] = `CIPHERTEXT_WIDTH'd4349168;
cipher_text[18] = `CIPHERTEXT_WIDTH'd14556581;
cipher_text[19] = `CIPHERTEXT_WIDTH'd8403081;
cipher_text[20] = `CIPHERTEXT_WIDTH'd15598499;
cipher_text[21] = `CIPHERTEXT_WIDTH'd13579739;
cipher_text[22] = `CIPHERTEXT_WIDTH'd7144212;
cipher_text[23] = `CIPHERTEXT_WIDTH'd13506946;
cipher_text[24] = `CIPHERTEXT_WIDTH'd8376866;
cipher_text[25] = `CIPHERTEXT_WIDTH'd2337756;
cipher_text[26] = `CIPHERTEXT_WIDTH'd4942005;
cipher_text[27] = `CIPHERTEXT_WIDTH'd5804784;
cipher_text[28] = `CIPHERTEXT_WIDTH'd13437089;
cipher_text[29] = `CIPHERTEXT_WIDTH'd8277705;
cipher_text[30] = `CIPHERTEXT_WIDTH'd15694784;
cipher_text[31] = `CIPHERTEXT_WIDTH'd6151379;
cipher_text[32] = `CIPHERTEXT_WIDTH'd1971770;
cipher_text[33] = `CIPHERTEXT_WIDTH'd15952769;
cipher_text[34] = `CIPHERTEXT_WIDTH'd1499190;
cipher_text[35] = `CIPHERTEXT_WIDTH'd3412154;
cipher_text[36] = `CIPHERTEXT_WIDTH'd1047633;
cipher_text[37] = `CIPHERTEXT_WIDTH'd652569;
cipher_text[38] = `CIPHERTEXT_WIDTH'd3805657;
cipher_text[39] = `CIPHERTEXT_WIDTH'd9098109;
cipher_text[40] = `CIPHERTEXT_WIDTH'd16637157;
cipher_text[41] = `CIPHERTEXT_WIDTH'd2034663;
cipher_text[42] = `CIPHERTEXT_WIDTH'd16616050;
cipher_text[43] = `CIPHERTEXT_WIDTH'd9114304;
cipher_text[44] = `CIPHERTEXT_WIDTH'd9778488;
cipher_text[45] = `CIPHERTEXT_WIDTH'd9073376;
cipher_text[46] = `CIPHERTEXT_WIDTH'd10544590;
cipher_text[47] = `CIPHERTEXT_WIDTH'd11452727;
cipher_text[48] = `CIPHERTEXT_WIDTH'd10561725;
cipher_text[49] = `CIPHERTEXT_WIDTH'd10553321;
cipher_text[50] = `CIPHERTEXT_WIDTH'd2982148;
cipher_text[51] = `CIPHERTEXT_WIDTH'd11214587;
cipher_text[52] = `CIPHERTEXT_WIDTH'd13577215;
cipher_text[53] = `CIPHERTEXT_WIDTH'd13850796;
cipher_text[54] = `CIPHERTEXT_WIDTH'd1260398;
cipher_text[55] = `CIPHERTEXT_WIDTH'd7999912;
cipher_text[56] = `CIPHERTEXT_WIDTH'd9146479;
cipher_text[57] = `CIPHERTEXT_WIDTH'd1675497;
cipher_text[58] = `CIPHERTEXT_WIDTH'd3817663;
cipher_text[59] = `CIPHERTEXT_WIDTH'd1917521;
cipher_text[60] = `CIPHERTEXT_WIDTH'd2407529;
cipher_text[61] = `CIPHERTEXT_WIDTH'd174226;
cipher_text[62] = `CIPHERTEXT_WIDTH'd2260261;
cipher_text[63] = `CIPHERTEXT_WIDTH'd13397535;
cipher_text[64] = `CIPHERTEXT_WIDTH'd4467971;
cipher_text[65] = `CIPHERTEXT_WIDTH'd8868997;
cipher_text[66] = `CIPHERTEXT_WIDTH'd12732193;
cipher_text[67] = `CIPHERTEXT_WIDTH'd13481853;
cipher_text[68] = `CIPHERTEXT_WIDTH'd9510872;
cipher_text[69] = `CIPHERTEXT_WIDTH'd14060507;
cipher_text[70] = `CIPHERTEXT_WIDTH'd3386842;
cipher_text[71] = `CIPHERTEXT_WIDTH'd11759078;
cipher_text[72] = `CIPHERTEXT_WIDTH'd337876;
cipher_text[73] = `CIPHERTEXT_WIDTH'd2850441;
cipher_text[74] = `CIPHERTEXT_WIDTH'd67473;
cipher_text[75] = `CIPHERTEXT_WIDTH'd388354;
cipher_text[76] = `CIPHERTEXT_WIDTH'd12768149;
cipher_text[77] = `CIPHERTEXT_WIDTH'd13135223;
cipher_text[78] = `CIPHERTEXT_WIDTH'd11699177;
cipher_text[79] = `CIPHERTEXT_WIDTH'd11051305;
cipher_text[80] = `CIPHERTEXT_WIDTH'd7192398;
cipher_text[81] = `CIPHERTEXT_WIDTH'd2619412;
cipher_text[82] = `CIPHERTEXT_WIDTH'd5327247;
cipher_text[83] = `CIPHERTEXT_WIDTH'd5545679;
cipher_text[84] = `CIPHERTEXT_WIDTH'd8382325;
cipher_text[85] = `CIPHERTEXT_WIDTH'd4552728;
cipher_text[86] = `CIPHERTEXT_WIDTH'd11571413;
cipher_text[87] = `CIPHERTEXT_WIDTH'd5855897;
cipher_text[88] = `CIPHERTEXT_WIDTH'd703609;
cipher_text[89] = `CIPHERTEXT_WIDTH'd8902068;
cipher_text[90] = `CIPHERTEXT_WIDTH'd7196819;
cipher_text[91] = `CIPHERTEXT_WIDTH'd3384420;
cipher_text[92] = `CIPHERTEXT_WIDTH'd619998;
cipher_text[93] = `CIPHERTEXT_WIDTH'd11533546;
cipher_text[94] = `CIPHERTEXT_WIDTH'd5191834;
cipher_text[95] = `CIPHERTEXT_WIDTH'd15203138;
cipher_text[96] = `CIPHERTEXT_WIDTH'd513796;
cipher_text[97] = `CIPHERTEXT_WIDTH'd8558688;
cipher_text[98] = `CIPHERTEXT_WIDTH'd14235763;
cipher_text[99] = `CIPHERTEXT_WIDTH'd6109758;
cipher_text[100] = `CIPHERTEXT_WIDTH'd9182325;
cipher_text[101] = `CIPHERTEXT_WIDTH'd14300425;
cipher_text[102] = `CIPHERTEXT_WIDTH'd15400992;
cipher_text[103] = `CIPHERTEXT_WIDTH'd12053924;
cipher_text[104] = `CIPHERTEXT_WIDTH'd9135234;
cipher_text[105] = `CIPHERTEXT_WIDTH'd9422654;
cipher_text[106] = `CIPHERTEXT_WIDTH'd7333683;
cipher_text[107] = `CIPHERTEXT_WIDTH'd14486643;
cipher_text[108] = `CIPHERTEXT_WIDTH'd513838;
cipher_text[109] = `CIPHERTEXT_WIDTH'd11264730;
cipher_text[110] = `CIPHERTEXT_WIDTH'd16671020;
cipher_text[111] = `CIPHERTEXT_WIDTH'd1057693;
cipher_text[112] = `CIPHERTEXT_WIDTH'd10342734;
cipher_text[113] = `CIPHERTEXT_WIDTH'd4345352;
cipher_text[114] = `CIPHERTEXT_WIDTH'd10962983;
cipher_text[115] = `CIPHERTEXT_WIDTH'd15959559;
cipher_text[116] = `CIPHERTEXT_WIDTH'd5152897;
cipher_text[117] = `CIPHERTEXT_WIDTH'd11017920;
cipher_text[118] = `CIPHERTEXT_WIDTH'd9316744;
cipher_text[119] = `CIPHERTEXT_WIDTH'd16277093;
cipher_text[120] = `CIPHERTEXT_WIDTH'd5700283;
cipher_text[121] = `CIPHERTEXT_WIDTH'd3948264;
cipher_text[122] = `CIPHERTEXT_WIDTH'd10658709;
cipher_text[123] = `CIPHERTEXT_WIDTH'd6705083;
cipher_text[124] = `CIPHERTEXT_WIDTH'd6624667;
cipher_text[125] = `CIPHERTEXT_WIDTH'd9678162;
cipher_text[126] = `CIPHERTEXT_WIDTH'd476819;
cipher_text[127] = `CIPHERTEXT_WIDTH'd411030;
cipher_text[128] = `CIPHERTEXT_WIDTH'd7934873;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
row = 128;
skentry = secret_key[128];
ctentry = cipher_text[128];
#20;
$display("Result = %d", result); assert(result == expected);

$finish;
end
endmodule