../results/user_proj_example.lef