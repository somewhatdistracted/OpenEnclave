module sram
#(
    parameter DATA_WIDTH = 32,
    parameter ADDR_WIDTH = 10,
    parameter DEPTH = 1024
)
(
    input clk,

    input in_wen,
    input [ADDR_WIDTH - 1 : 0] in_wadr,
    input [DATA_WIDTH - 1 : 0] in_wdata,

    input out_wen,
    input [ADDR_WIDTH - 1 : 0] out_wadr,
    input [DATA_WIDTH - 1 : 0] out_wdata,

    input op1_ren,
    input [ADDR_WIDTH - 1 : 0] op1_radr,
    output [DATA_WIDTH - 1 : 0] op1_rdata,

    input op2_ren,
    input [ADDR_WIDTH - 1 : 0] op2_radr,
    output [DATA_WIDTH - 1 : 0] op2_rdata,
    
    input out_ren,
    input [ADDR_WIDTH - 1 : 0] out_radr,
    output [DATA_WIDTH - 1 : 0] out_rdata
);

    genvar x, y;
    generate
        wire [DATA_WIDTH - 1 : 0] op1_rdata_w [DEPTH/256 - 1 : 0]; 
        reg  [ADDR_WIDTH - 1 : 0] op1_radr_r;
        wire [DATA_WIDTH - 1 : 0] op2_rdata_w [DEPTH/256 - 1 : 0]; 
        reg  [ADDR_WIDTH - 1 : 0] op2_radr_r;
        wire [DATA_WIDTH - 1 : 0] out_rdata_w [DEPTH/256 - 1 : 0]; 
        reg  [ADDR_WIDTH - 1 : 0] out_radr_r;

        always @ (posedge clk) begin
            op1_radr_r <= op1_radr;
            op2_radr_r <= op2_radr;
            out_radr_r <= out_radr;
        end 

        // op1
        for (x = 0; x < DATA_WIDTH/32; x = x + 1) begin: width_macro1
            for (y = 0; y < DEPTH/256; y = y + 1) begin: depth_macro1
                // note: Excerpted from EE272 Sram Wrapper:
                // note: The default behavioral model generated by OpenRAM has an arbitrary
                //       delay of 3ns. Since the SRAM data is only valid for half a cycle
                //       any delay < half a cycle will not affect the simulation result.
                //       Since we will try to push for a clock period of 5ns, we manually
                //       changed the delay number to 1ns (< 2.5ns) to prevent functional error.
                sky130_sram_1kbyte_1rw1r_32x256_8 sram1 (
                    .clk0(clk),
                    .csb0(~(in_wen && (in_wadr[ADDR_WIDTH - 1 : 8] == y))),
                    .web0(~(in_wen && (in_wadr[ADDR_WIDTH - 1 : 8] == y))), // And wadr in range
                    .wmask0(4'hF),
                    .addr0(in_wadr[7:0]),
                    .din0(in_wdata[32*(x+1)-1 : 32*x]),
                    .dout0(),
                    .clk1(clk),
                    .csb1(~(op1_ren && (op1_radr[ADDR_WIDTH - 1 : 8] == y))), // And radr in range
                    .addr1(op1_radr[7:0]),
                    .dout1(op1_rdata_w[y][32*(x+1)-1 : 32*x])
                );
            end
        end

        // op2
        for (x = 0; x < DATA_WIDTH/32; x = x + 1) begin: width_macro2
            for (y = 0; y < DEPTH/256; y = y + 1) begin: depth_macro2
                // note: Excerpted from EE272 Sram Wrapper:
                // note: The default behavioral model generated by OpenRAM has an arbitrary
                //       delay of 3ns. Since the SRAM data is only valid for half a cycle
                //       any delay < half a cycle will not affect the simulation result.
                //       Since we will try to push for a clock period of 5ns, we manually
                //       changed the delay number to 1ns (< 2.5ns) to prevent functional error.
                sky130_sram_1kbyte_1rw1r_32x256_8 sram2 (
                    .clk0(clk),
                    .csb0(~(in_wen && (in_wadr[ADDR_WIDTH - 1 : 8] == y))),
                    .web0(~(in_wen && (in_wadr[ADDR_WIDTH - 1 : 8] == y))), // And wadr in range
                    .wmask0(4'hF),
                    .addr0(in_wadr[7:0]),
                    .din0(in_wdata[32*(x+1)-1 : 32*x]),
                    .dout0(),
                    .clk1(clk),
                    .csb1(~(op2_ren && (op2_radr[ADDR_WIDTH - 1 : 8] == y))), // And radr in range
                    .addr1(op2_radr[7:0]),
                    .dout1(op2_rdata_w[y][32*(x+1)-1 : 32*x])
                );
            end
        end

        // out
        for (x = 0; x < DATA_WIDTH/32; x = x + 1) begin: width_macro3
            for (y = 0; y < DEPTH/256; y = y + 1) begin: depth_macro3
                // note: Excerpted from EE272 Sram Wrapper:
                // note: The default behavioral model generated by OpenRAM has an arbitrary
                //       delay of 3ns. Since the SRAM data is only valid for half a cycle
                //       any delay < half a cycle will not affect the simulation result.
                //       Since we will try to push for a clock period of 5ns, we manually
                //       changed the delay number to 1ns (< 2.5ns) to prevent functional error.
                sky130_sram_1kbyte_1rw1r_32x256_8 sram3 (
                    .clk0(clk),
                    .csb0(~(out_wen && (out_wadr[ADDR_WIDTH - 1 : 8] == y))),
                    .web0(~(out_wen && (out_wadr[ADDR_WIDTH - 1 : 8] == y))), // And wadr in range
                    .wmask0(4'hF),
                    .addr0(out_wadr[7:0]),
                    .din0(out_wdata[32*(x+1)-1 : 32*x]),
                    .dout0(),
                    .clk1(clk),
                    .csb1(~(out_ren && (out_radr[ADDR_WIDTH - 1 : 8] == y))), // And radr in range
                    .addr1(out_radr[7:0]),
                    .dout1(out_rdata_w[y][32*(x+1)-1 : 32*x])
                );
            end
        end

    endgenerate

    assign op1_rdata = op1_rdata_w[op1_radr_r[ADDR_WIDTH - 1 : 8]];
    assign op2_rdata = op2_rdata_w[op2_radr_r[ADDR_WIDTH - 1 : 8]];
    assign out_rdata = out_rdata_w[out_radr_r[ADDR_WIDTH - 1 : 8]];

endmodule
