/home/users/ianpmac/EE372-Project/skywater-digital-flow/HEModules/build/5-skywater-130nm/view-standard/stdcells.lef