`define PLAINTEXT_MODULUS 32
`define PLAINTEXT_WIDTH 5
`define DIMENSION 128
`define CIPHERTEXT_MODULUS 16777216
`define CIPHERTEXT_WIDTH 24
`define BIG_N 6425

module homomorphic_multiply_tb;

    reg clk;
    reg rst_n;
    reg signed [`CIPHERTEXT_WIDTH-1:0] ciphertext_entry;
    reg [`DIMENSION:0] row;
    reg ciphertext_select;
    reg en;
    wire signed [`CIPHERTEXT_WIDTH-1:0] result;
    reg signed [`CIPHERTEXT_WIDTH-1:0] expected;

    always #10 clk = ~clk;

    homomorphic_multiply #(
        .PLAINTEXT_MODULUS(`PLAINTEXT_MODULUS),
        .PLAINTEXT_WIDTH(`PLAINTEXT_WIDTH),
        .CIPHERTEXT_MODULUS(`CIPHERTEXT_MODULUS),
        .CIPHERTEXT_WIDTH(`CIPHERTEXT_WIDTH),
        .DIMENSION(`DIMENSION),
        .BIG_N(`BIG_N)
    ) homomorphic_inst (
        .clk(clk),
        .rst_n(rst_n),
        .ciphertext_entry(ciphertext_entry),
        .row(row),
        .ciphertext_select(ciphertext_select),
        .en(en),
        .result_partial(result)
    );

    initial begin
        clk = 0;
        ciphertext_select = 0;
        row = 0;
        ciphertext_entry = 0;

en=0;
rst_n=0;
#100;
rst_n=1;
#100;
en=1;
#20;
ciphertext_select = 0;
row = 0;
ciphertext_entry =4120072;
#20;
row = 1;
ciphertext_entry =6284281;
#20;
row = 2;
ciphertext_entry =9554369;
#20;
row = 3;
ciphertext_entry =9222648;
#20;
row = 4;
ciphertext_entry =14029513;
#20;
row = 5;
ciphertext_entry =920679;
#20;
row = 6;
ciphertext_entry =6769264;
#20;
row = 7;
ciphertext_entry =6205512;
#20;
row = 8;
ciphertext_entry =1773446;
#20;
row = 9;
ciphertext_entry =6684276;
#20;
row = 10;
ciphertext_entry =9722837;
#20;
row = 11;
ciphertext_entry =4321959;
#20;
row = 12;
ciphertext_entry =11817387;
#20;
row = 13;
ciphertext_entry =5563913;
#20;
row = 14;
ciphertext_entry =3723396;
#20;
row = 15;
ciphertext_entry =8439575;
#20;
row = 16;
ciphertext_entry =14213459;
#20;
row = 17;
ciphertext_entry =5560018;
#20;
row = 18;
ciphertext_entry =16574204;
#20;
row = 19;
ciphertext_entry =2393083;
#20;
row = 20;
ciphertext_entry =819119;
#20;
row = 21;
ciphertext_entry =1197976;
#20;
row = 22;
ciphertext_entry =12235107;
#20;
row = 23;
ciphertext_entry =5764253;
#20;
row = 24;
ciphertext_entry =8257962;
#20;
row = 25;
ciphertext_entry =4156060;
#20;
row = 26;
ciphertext_entry =8273660;
#20;
row = 27;
ciphertext_entry =3700265;
#20;
row = 28;
ciphertext_entry =407900;
#20;
row = 29;
ciphertext_entry =14935934;
#20;
row = 30;
ciphertext_entry =16684946;
#20;
row = 31;
ciphertext_entry =6576630;
#20;
row = 32;
ciphertext_entry =16224260;
#20;
row = 33;
ciphertext_entry =13312306;
#20;
row = 34;
ciphertext_entry =12308926;
#20;
row = 35;
ciphertext_entry =1609843;
#20;
row = 36;
ciphertext_entry =7681394;
#20;
row = 37;
ciphertext_entry =11721859;
#20;
row = 38;
ciphertext_entry =1166532;
#20;
row = 39;
ciphertext_entry =910729;
#20;
row = 40;
ciphertext_entry =3295280;
#20;
row = 41;
ciphertext_entry =12641252;
#20;
row = 42;
ciphertext_entry =4629394;
#20;
row = 43;
ciphertext_entry =4699428;
#20;
row = 44;
ciphertext_entry =8710274;
#20;
row = 45;
ciphertext_entry =8520077;
#20;
row = 46;
ciphertext_entry =8454874;
#20;
row = 47;
ciphertext_entry =3193917;
#20;
row = 48;
ciphertext_entry =15758932;
#20;
row = 49;
ciphertext_entry =3292319;
#20;
row = 50;
ciphertext_entry =12173657;
#20;
row = 51;
ciphertext_entry =10776473;
#20;
row = 52;
ciphertext_entry =11208448;
#20;
row = 53;
ciphertext_entry =6958343;
#20;
row = 54;
ciphertext_entry =2211680;
#20;
row = 55;
ciphertext_entry =15302981;
#20;
row = 56;
ciphertext_entry =8066182;
#20;
row = 57;
ciphertext_entry =9530345;
#20;
row = 58;
ciphertext_entry =15757222;
#20;
row = 59;
ciphertext_entry =7360780;
#20;
row = 60;
ciphertext_entry =6934056;
#20;
row = 61;
ciphertext_entry =13002921;
#20;
row = 62;
ciphertext_entry =12890229;
#20;
row = 63;
ciphertext_entry =12604482;
#20;
row = 64;
ciphertext_entry =13966699;
#20;
row = 65;
ciphertext_entry =8475669;
#20;
row = 66;
ciphertext_entry =6259879;
#20;
row = 67;
ciphertext_entry =2836796;
#20;
row = 68;
ciphertext_entry =6454473;
#20;
row = 69;
ciphertext_entry =2966774;
#20;
row = 70;
ciphertext_entry =9322038;
#20;
row = 71;
ciphertext_entry =8610819;
#20;
row = 72;
ciphertext_entry =3982302;
#20;
row = 73;
ciphertext_entry =3599882;
#20;
row = 74;
ciphertext_entry =16129971;
#20;
row = 75;
ciphertext_entry =15768454;
#20;
row = 76;
ciphertext_entry =4668831;
#20;
row = 77;
ciphertext_entry =12705696;
#20;
row = 78;
ciphertext_entry =13550561;
#20;
row = 79;
ciphertext_entry =5882296;
#20;
row = 80;
ciphertext_entry =4599916;
#20;
row = 81;
ciphertext_entry =2997892;
#20;
row = 82;
ciphertext_entry =527561;
#20;
row = 83;
ciphertext_entry =15849075;
#20;
row = 84;
ciphertext_entry =14035033;
#20;
row = 85;
ciphertext_entry =179944;
#20;
row = 86;
ciphertext_entry =6025078;
#20;
row = 87;
ciphertext_entry =5841670;
#20;
row = 88;
ciphertext_entry =1944946;
#20;
row = 89;
ciphertext_entry =11061664;
#20;
row = 90;
ciphertext_entry =8002903;
#20;
row = 91;
ciphertext_entry =13503603;
#20;
row = 92;
ciphertext_entry =4650609;
#20;
row = 93;
ciphertext_entry =7016761;
#20;
row = 94;
ciphertext_entry =9994392;
#20;
row = 95;
ciphertext_entry =4469116;
#20;
row = 96;
ciphertext_entry =10251515;
#20;
row = 97;
ciphertext_entry =1324426;
#20;
row = 98;
ciphertext_entry =7465021;
#20;
row = 99;
ciphertext_entry =7027450;
#20;
row = 100;
ciphertext_entry =2059977;
#20;
row = 101;
ciphertext_entry =9487252;
#20;
row = 102;
ciphertext_entry =14515492;
#20;
row = 103;
ciphertext_entry =7740267;
#20;
row = 104;
ciphertext_entry =9114581;
#20;
row = 105;
ciphertext_entry =4082121;
#20;
row = 106;
ciphertext_entry =7933236;
#20;
row = 107;
ciphertext_entry =11318175;
#20;
row = 108;
ciphertext_entry =9992298;
#20;
row = 109;
ciphertext_entry =1521440;
#20;
row = 110;
ciphertext_entry =3433450;
#20;
row = 111;
ciphertext_entry =10860466;
#20;
row = 112;
ciphertext_entry =12703542;
#20;
row = 113;
ciphertext_entry =8774313;
#20;
row = 114;
ciphertext_entry =3337481;
#20;
row = 115;
ciphertext_entry =12574408;
#20;
row = 116;
ciphertext_entry =14061099;
#20;
row = 117;
ciphertext_entry =1439866;
#20;
row = 118;
ciphertext_entry =14967150;
#20;
row = 119;
ciphertext_entry =9507671;
#20;
row = 120;
ciphertext_entry =6631663;
#20;
row = 121;
ciphertext_entry =2978676;
#20;
row = 122;
ciphertext_entry =6323747;
#20;
row = 123;
ciphertext_entry =9977585;
#20;
row = 124;
ciphertext_entry =1436668;
#20;
row = 125;
ciphertext_entry =15070764;
#20;
row = 126;
ciphertext_entry =16717579;
#20;
row = 127;
ciphertext_entry =15542931;
#20;
row = 128;
ciphertext_entry =1757079;
#20;
ciphertext_select = 1;
row = 0;
ciphertext_entry =4120072;
#20;
$display("Result = %d", result); assert(result ==9923152);
row = 1;
ciphertext_entry =6284281;
#20;
$display("Result = %d", result); assert(result ==10604114);
row = 2;
ciphertext_entry =9554369;
#20;
$display("Result = %d", result); assert(result ==10624501);
row = 3;
ciphertext_entry =9222648;
#20;
$display("Result = %d", result); assert(result ==11457768);
row = 4;
ciphertext_entry =14029513;
#20;
$display("Result = %d", result); assert(result ==9802779);
row = 5;
ciphertext_entry =920679;
#20;
$display("Result = %d", result); assert(result ==14849560);
row = 6;
ciphertext_entry =6769264;
#20;
$display("Result = %d", result); assert(result ==5358250);
row = 7;
ciphertext_entry =6205512;
#20;
$display("Result = %d", result); assert(result ==13910290);
row = 8;
ciphertext_entry =1773446;
#20;
$display("Result = %d", result); assert(result ==2442549);
row = 9;
ciphertext_entry =6684276;
#20;
$display("Result = %d", result); assert(result ==347780);
row = 10;
ciphertext_entry =9722837;
#20;
$display("Result = %d", result); assert(result ==5467550);
row = 11;
ciphertext_entry =4321959;
#20;
$display("Result = %d", result); assert(result ==6281473);
row = 12;
ciphertext_entry =11817387;
#20;
$display("Result = %d", result); assert(result ==13317112);
row = 13;
ciphertext_entry =5563913;
#20;
$display("Result = %d", result); assert(result ==6240175);
row = 14;
ciphertext_entry =3723396;
#20;
$display("Result = %d", result); assert(result ==15338147);
row = 15;
ciphertext_entry =8439575;
#20;
$display("Result = %d", result); assert(result ==1561049);
row = 16;
ciphertext_entry =14213459;
#20;
$display("Result = %d", result); assert(result ==15344975);
row = 17;
ciphertext_entry =5560018;
#20;
$display("Result = %d", result); assert(result ==758843);
row = 18;
ciphertext_entry =16574204;
#20;
$display("Result = %d", result); assert(result ==1595245);
row = 19;
ciphertext_entry =2393083;
#20;
$display("Result = %d", result); assert(result ==12169173);
row = 20;
ciphertext_entry =819119;
#20;
$display("Result = %d", result); assert(result ==357138);
row = 21;
ciphertext_entry =1197976;
#20;
$display("Result = %d", result); assert(result ==9503935);
row = 22;
ciphertext_entry =12235107;
#20;
$display("Result = %d", result); assert(result ==14255452);
row = 23;
ciphertext_entry =5764253;
#20;
$display("Result = %d", result); assert(result ==12895925);
row = 24;
ciphertext_entry =8257962;
#20;
$display("Result = %d", result); assert(result ==12208066);
row = 25;
ciphertext_entry =4156060;
#20;
$display("Result = %d", result); assert(result ==1936401);
row = 26;
ciphertext_entry =8273660;
#20;
$display("Result = %d", result); assert(result ==2242229);
row = 27;
ciphertext_entry =3700265;
#20;
$display("Result = %d", result); assert(result ==12319695);
row = 28;
ciphertext_entry =407900;
#20;
$display("Result = %d", result); assert(result ==14385287);
row = 29;
ciphertext_entry =14935934;
#20;
$display("Result = %d", result); assert(result ==2041031);
row = 30;
ciphertext_entry =16684946;
#20;
$display("Result = %d", result); assert(result ==4896781);
row = 31;
ciphertext_entry =6576630;
#20;
$display("Result = %d", result); assert(result ==13067545);
row = 32;
ciphertext_entry =16224260;
#20;
$display("Result = %d", result); assert(result ==13153511);
row = 33;
ciphertext_entry =13312306;
#20;
$display("Result = %d", result); assert(result ==9910059);
row = 34;
ciphertext_entry =12308926;
#20;
$display("Result = %d", result); assert(result ==7533426);
row = 35;
ciphertext_entry =1609843;
#20;
$display("Result = %d", result); assert(result ==3998290);
row = 36;
ciphertext_entry =7681394;
#20;
$display("Result = %d", result); assert(result ==2193572);
row = 37;
ciphertext_entry =11721859;
#20;
$display("Result = %d", result); assert(result ==8024581);
row = 38;
ciphertext_entry =1166532;
#20;
$display("Result = %d", result); assert(result ==4495659);
row = 39;
ciphertext_entry =910729;
#20;
$display("Result = %d", result); assert(result ==9879486);
row = 40;
ciphertext_entry =3295280;
#20;
$display("Result = %d", result); assert(result ==8574680);
row = 41;
ciphertext_entry =12641252;
#20;
$display("Result = %d", result); assert(result ==4211031);
row = 42;
ciphertext_entry =4629394;
#20;
$display("Result = %d", result); assert(result ==12432166);
row = 43;
ciphertext_entry =4699428;
#20;
$display("Result = %d", result); assert(result ==2496192);
row = 44;
ciphertext_entry =8710274;
#20;
$display("Result = %d", result); assert(result ==12299255);
row = 45;
ciphertext_entry =8520077;
#20;
$display("Result = %d", result); assert(result ==6715150);
row = 46;
ciphertext_entry =8454874;
#20;
$display("Result = %d", result); assert(result ==4252658);
row = 47;
ciphertext_entry =3193917;
#20;
$display("Result = %d", result); assert(result ==6934477);
row = 48;
ciphertext_entry =15758932;
#20;
$display("Result = %d", result); assert(result ==16750453);
row = 49;
ciphertext_entry =3292319;
#20;
$display("Result = %d", result); assert(result ==3525942);
row = 50;
ciphertext_entry =12173657;
#20;
$display("Result = %d", result); assert(result ==15640798);
row = 51;
ciphertext_entry =10776473;
#20;
$display("Result = %d", result); assert(result ==15469787);
row = 52;
ciphertext_entry =11208448;
#20;
$display("Result = %d", result); assert(result ==4138793);
row = 53;
ciphertext_entry =6958343;
#20;
$display("Result = %d", result); assert(result ==9606170);
row = 54;
ciphertext_entry =2211680;
#20;
$display("Result = %d", result); assert(result ==4808192);
row = 55;
ciphertext_entry =15302981;
#20;
$display("Result = %d", result); assert(result ==3144266);
row = 56;
ciphertext_entry =8066182;
#20;
$display("Result = %d", result); assert(result ==13849080);
row = 57;
ciphertext_entry =9530345;
#20;
$display("Result = %d", result); assert(result ==1049850);
row = 58;
ciphertext_entry =15757222;
#20;
$display("Result = %d", result); assert(result ==14725264);
row = 59;
ciphertext_entry =7360780;
#20;
$display("Result = %d", result); assert(result ==16442460);
row = 60;
ciphertext_entry =6934056;
#20;
$display("Result = %d", result); assert(result ==9653656);
row = 61;
ciphertext_entry =13002921;
#20;
$display("Result = %d", result); assert(result ==4257264);
row = 62;
ciphertext_entry =12890229;
#20;
$display("Result = %d", result); assert(result ==6662747);
row = 63;
ciphertext_entry =12604482;
#20;
$display("Result = %d", result); assert(result ==5202101);
row = 64;
ciphertext_entry =13966699;
#20;
$display("Result = %d", result); assert(result ==835633);
row = 65;
ciphertext_entry =8475669;
#20;
$display("Result = %d", result); assert(result ==8718407);
row = 66;
ciphertext_entry =6259879;
#20;
$display("Result = %d", result); assert(result ==9225502);
row = 67;
ciphertext_entry =2836796;
#20;
$display("Result = %d", result); assert(result ==12328006);
row = 68;
ciphertext_entry =6454473;
#20;
$display("Result = %d", result); assert(result ==8530830);
row = 69;
ciphertext_entry =2966774;
#20;
$display("Result = %d", result); assert(result ==2437740);
row = 70;
ciphertext_entry =9322038;
#20;
$display("Result = %d", result); assert(result ==12334375);
row = 71;
ciphertext_entry =8610819;
#20;
$display("Result = %d", result); assert(result ==5241277);
row = 72;
ciphertext_entry =3982302;
#20;
$display("Result = %d", result); assert(result ==16362660);
row = 73;
ciphertext_entry =3599882;
#20;
$display("Result = %d", result); assert(result ==6779140);
row = 74;
ciphertext_entry =16129971;
#20;
$display("Result = %d", result); assert(result ==514626);
row = 75;
ciphertext_entry =15768454;
#20;
$display("Result = %d", result); assert(result ==5567534);
row = 76;
ciphertext_entry =4668831;
#20;
$display("Result = %d", result); assert(result ==6367087);
row = 77;
ciphertext_entry =12705696;
#20;
$display("Result = %d", result); assert(result ==12717531);
row = 78;
ciphertext_entry =13550561;
#20;
$display("Result = %d", result); assert(result ==12915171);
row = 79;
ciphertext_entry =5882296;
#20;
$display("Result = %d", result); assert(result ==2079772);
row = 80;
ciphertext_entry =4599916;
#20;
$display("Result = %d", result); assert(result ==5795499);
row = 81;
ciphertext_entry =2997892;
#20;
$display("Result = %d", result); assert(result ==9228725);
row = 82;
ciphertext_entry =527561;
#20;
$display("Result = %d", result); assert(result ==15565651);
row = 83;
ciphertext_entry =15849075;
#20;
$display("Result = %d", result); assert(result ==7266952);
row = 84;
ciphertext_entry =14035033;
#20;
$display("Result = %d", result); assert(result ==15860414);
row = 85;
ciphertext_entry =179944;
#20;
$display("Result = %d", result); assert(result ==10752462);
row = 86;
ciphertext_entry =6025078;
#20;
$display("Result = %d", result); assert(result ==13900413);
row = 87;
ciphertext_entry =5841670;
#20;
$display("Result = %d", result); assert(result ==15635283);
row = 88;
ciphertext_entry =1944946;
#20;
$display("Result = %d", result); assert(result ==16670734);
row = 89;
ciphertext_entry =11061664;
#20;
$display("Result = %d", result); assert(result ==4872224);
row = 90;
ciphertext_entry =8002903;
#20;
$display("Result = %d", result); assert(result ==16203638);
row = 91;
ciphertext_entry =13503603;
#20;
$display("Result = %d", result); assert(result ==15689296);
row = 92;
ciphertext_entry =4650609;
#20;
$display("Result = %d", result); assert(result ==12970492);
row = 93;
ciphertext_entry =7016761;
#20;
$display("Result = %d", result); assert(result ==8034441);
row = 94;
ciphertext_entry =9994392;
#20;
$display("Result = %d", result); assert(result ==11661944);
row = 95;
ciphertext_entry =4469116;
#20;
$display("Result = %d", result); assert(result ==10385303);
row = 96;
ciphertext_entry =10251515;
#20;
$display("Result = %d", result); assert(result ==13232846);
row = 97;
ciphertext_entry =1324426;
#20;
$display("Result = %d", result); assert(result ==1068183);
row = 98;
ciphertext_entry =7465021;
#20;
$display("Result = %d", result); assert(result ==5368340);
row = 99;
ciphertext_entry =7027450;
#20;
$display("Result = %d", result); assert(result ==4956761);
row = 100;
ciphertext_entry =2059977;
#20;
$display("Result = %d", result); assert(result ==7973119);
row = 101;
ciphertext_entry =9487252;
#20;
$display("Result = %d", result); assert(result ==8674871);
row = 102;
ciphertext_entry =14515492;
#20;
$display("Result = %d", result); assert(result ==9671497);
row = 103;
ciphertext_entry =7740267;
#20;
$display("Result = %d", result); assert(result ==12101602);
row = 104;
ciphertext_entry =9114581;
#20;
$display("Result = %d", result); assert(result ==10691137);
row = 105;
ciphertext_entry =4082121;
#20;
$display("Result = %d", result); assert(result ==11246931);
row = 106;
ciphertext_entry =7933236;
#20;
$display("Result = %d", result); assert(result ==12435017);
row = 107;
ciphertext_entry =11318175;
#20;
$display("Result = %d", result); assert(result ==2775339);
row = 108;
ciphertext_entry =9992298;
#20;
$display("Result = %d", result); assert(result ==1745858);
row = 109;
ciphertext_entry =1521440;
#20;
$display("Result = %d", result); assert(result ==9098908);
row = 110;
ciphertext_entry =3433450;
#20;
$display("Result = %d", result); assert(result ==213851);
row = 111;
ciphertext_entry =10860466;
#20;
$display("Result = %d", result); assert(result ==7204705);
row = 112;
ciphertext_entry =12703542;
#20;
$display("Result = %d", result); assert(result ==1866787);
row = 113;
ciphertext_entry =8774313;
#20;
$display("Result = %d", result); assert(result ==7436481);
row = 114;
ciphertext_entry =3337481;
#20;
$display("Result = %d", result); assert(result ==10024552);
row = 115;
ciphertext_entry =12574408;
#20;
$display("Result = %d", result); assert(result ==9358787);
row = 116;
ciphertext_entry =14061099;
#20;
$display("Result = %d", result); assert(result ==9189172);
row = 117;
ciphertext_entry =1439866;
#20;
$display("Result = %d", result); assert(result ==3999764);
row = 118;
ciphertext_entry =14967150;
#20;
$display("Result = %d", result); assert(result ==4923336);
row = 119;
ciphertext_entry =9507671;
#20;
$display("Result = %d", result); assert(result ==9061904);
row = 120;
ciphertext_entry =6631663;
#20;
$display("Result = %d", result); assert(result ==14975456);
row = 121;
ciphertext_entry =2978676;
#20;
$display("Result = %d", result); assert(result ==16580442);
row = 122;
ciphertext_entry =6323747;
#20;
$display("Result = %d", result); assert(result ==10838382);
row = 123;
ciphertext_entry =9977585;
#20;
$display("Result = %d", result); assert(result ==5925332);
row = 124;
ciphertext_entry =1436668;
#20;
$display("Result = %d", result); assert(result ==1484295);
row = 125;
ciphertext_entry =15070764;
#20;
$display("Result = %d", result); assert(result ==2879922);
row = 126;
ciphertext_entry =16717579;
#20;
$display("Result = %d", result); assert(result ==13496764);
row = 127;
ciphertext_entry =15542931;
#20;
$display("Result = %d", result); assert(result ==1125098);
row = 128;
ciphertext_entry =1757079;
#20;
$display("Result = %d", result); assert(result ==1686600);
ciphertext_select = 0;
row = 129;
#20;
$display("Result = %d", result); assert(result ==12943000);
row = 130;
#20;
$display("Result = %d", result); assert(result ==7184315);
row = 131;
#20;
$display("Result = %d", result); assert(result ==16709035);
row = 132;
#20;
$display("Result = %d", result); assert(result ==9437415);
row = 133;
#20;
$display("Result = %d", result); assert(result ==13624904);
row = 134;
#20;
$display("Result = %d", result); assert(result ==11718303);
row = 135;
#20;
$display("Result = %d", result); assert(result ==9597957);
row = 136;
#20;
$display("Result = %d", result); assert(result ==7347507);
row = 137;
#20;
$display("Result = %d", result); assert(result ==11208981);
row = 138;
#20;
$display("Result = %d", result); assert(result ==408655);
row = 139;
#20;
$display("Result = %d", result); assert(result ==9722872);
row = 140;
#20;
$display("Result = %d", result); assert(result ==16552882);
row = 141;
#20;
$display("Result = %d", result); assert(result ==13552504);
row = 142;
#20;
$display("Result = %d", result); assert(result ==12583643);
row = 143;
#20;
$display("Result = %d", result); assert(result ==5626295);
row = 144;
#20;
$display("Result = %d", result); assert(result ==4927822);
row = 145;
#20;
$display("Result = %d", result); assert(result ==8030070);
row = 146;
#20;
$display("Result = %d", result); assert(result ==6429037);
row = 147;
#20;
$display("Result = %d", result); assert(result ==7721948);
row = 148;
#20;
$display("Result = %d", result); assert(result ==15000260);
row = 149;
#20;
$display("Result = %d", result); assert(result ==1562785);
row = 150;
#20;
$display("Result = %d", result); assert(result ==13425433);
row = 151;
#20;
$display("Result = %d", result); assert(result ==14514716);
row = 152;
#20;
$display("Result = %d", result); assert(result ==15991241);
row = 153;
#20;
$display("Result = %d", result); assert(result ==1835818);
row = 154;
#20;
$display("Result = %d", result); assert(result ==3605338);
row = 155;
#20;
$display("Result = %d", result); assert(result ==9386371);
row = 156;
#20;
$display("Result = %d", result); assert(result ==268868);
row = 157;
#20;
$display("Result = %d", result); assert(result ==8625937);
row = 158;
#20;
$display("Result = %d", result); assert(result ==13187586);
row = 159;
#20;
$display("Result = %d", result); assert(result ==5329409);
row = 160;
#20;
$display("Result = %d", result); assert(result ==14639724);
row = 161;
#20;
$display("Result = %d", result); assert(result ==2275026);
row = 162;
#20;
$display("Result = %d", result); assert(result ==2583238);
row = 163;
#20;
$display("Result = %d", result); assert(result ==5922868);
row = 164;
#20;
$display("Result = %d", result); assert(result ==6663183);
row = 165;
#20;
$display("Result = %d", result); assert(result ==15821333);
row = 166;
#20;
$display("Result = %d", result); assert(result ==15383007);
row = 167;
#20;
$display("Result = %d", result); assert(result ==4240889);
row = 168;
#20;
$display("Result = %d", result); assert(result ==9175877);
row = 169;
#20;
$display("Result = %d", result); assert(result ==8173933);
row = 170;
#20;
$display("Result = %d", result); assert(result ==4120515);
row = 171;
#20;
$display("Result = %d", result); assert(result ==7189099);
row = 172;
#20;
$display("Result = %d", result); assert(result ==4583144);
row = 173;
#20;
$display("Result = %d", result); assert(result ==13959515);
row = 174;
#20;
$display("Result = %d", result); assert(result ==16117598);
row = 175;
#20;
$display("Result = %d", result); assert(result ==13429046);
row = 176;
#20;
$display("Result = %d", result); assert(result ==5728970);
row = 177;
#20;
$display("Result = %d", result); assert(result ==7633343);
row = 178;
#20;
$display("Result = %d", result); assert(result ==176181);
row = 179;
#20;
$display("Result = %d", result); assert(result ==11075074);
row = 180;
#20;
$display("Result = %d", result); assert(result ==4747374);
row = 181;
#20;
$display("Result = %d", result); assert(result ==13631616);
row = 182;
#20;
$display("Result = %d", result); assert(result ==15538593);
row = 183;
#20;
$display("Result = %d", result); assert(result ==6085531);
row = 184;
#20;
$display("Result = %d", result); assert(result ==16752747);
row = 185;
#20;
$display("Result = %d", result); assert(result ==15211948);
row = 186;
#20;
$display("Result = %d", result); assert(result ==7674077);
row = 187;
#20;
$display("Result = %d", result); assert(result ==15670921);
row = 188;
#20;
$display("Result = %d", result); assert(result ==8521939);
row = 189;
#20;
$display("Result = %d", result); assert(result ==14689012);
row = 190;
#20;
$display("Result = %d", result); assert(result ==14082155);
row = 191;
#20;
$display("Result = %d", result); assert(result ==491125);
row = 192;
#20;
$display("Result = %d", result); assert(result ==11229565);
row = 193;
#20;
$display("Result = %d", result); assert(result ==7907414);
row = 194;
#20;
$display("Result = %d", result); assert(result ==1141863);
row = 195;
#20;
$display("Result = %d", result); assert(result ==7217990);
row = 196;
#20;
$display("Result = %d", result); assert(result ==10546140);
row = 197;
#20;
$display("Result = %d", result); assert(result ==6298281);
row = 198;
#20;
$display("Result = %d", result); assert(result ==13839904);
row = 199;
#20;
$display("Result = %d", result); assert(result ==7069696);
row = 200;
#20;
$display("Result = %d", result); assert(result ==6743797);
row = 201;
#20;
$display("Result = %d", result); assert(result ==11113156);
row = 202;
#20;
$display("Result = %d", result); assert(result ==2059019);
row = 203;
#20;
$display("Result = %d", result); assert(result ==11442096);
row = 204;
#20;
$display("Result = %d", result); assert(result ==4959070);
row = 205;
#20;
$display("Result = %d", result); assert(result ==11270811);
row = 206;
#20;
$display("Result = %d", result); assert(result ==13427909);
row = 207;
#20;
$display("Result = %d", result); assert(result ==12957431);
row = 208;
#20;
$display("Result = %d", result); assert(result ==13785570);
row = 209;
#20;
$display("Result = %d", result); assert(result ==14465421);
row = 210;
#20;
$display("Result = %d", result); assert(result ==1376122);
row = 211;
#20;
$display("Result = %d", result); assert(result ==15113990);
row = 212;
#20;
$display("Result = %d", result); assert(result ==6433303);
row = 213;
#20;
$display("Result = %d", result); assert(result ==12620107);
row = 214;
#20;
$display("Result = %d", result); assert(result ==9604886);
row = 215;
#20;
$display("Result = %d", result); assert(result ==14581611);
row = 216;
#20;
$display("Result = %d", result); assert(result ==14960920);
row = 217;
#20;
$display("Result = %d", result); assert(result ==14705206);
row = 218;
#20;
$display("Result = %d", result); assert(result ==3177853);
row = 219;
#20;
$display("Result = %d", result); assert(result ==1977942);
row = 220;
#20;
$display("Result = %d", result); assert(result ==8954687);
row = 221;
#20;
$display("Result = %d", result); assert(result ==7194010);
row = 222;
#20;
$display("Result = %d", result); assert(result ==6651494);
row = 223;
#20;
$display("Result = %d", result); assert(result ==11825206);
row = 224;
#20;
$display("Result = %d", result); assert(result ==7492919);
row = 225;
#20;
$display("Result = %d", result); assert(result ==832218);
row = 226;
#20;
$display("Result = %d", result); assert(result ==16543572);
row = 227;
#20;
$display("Result = %d", result); assert(result ==16422044);
row = 228;
#20;
$display("Result = %d", result); assert(result ==4998587);
row = 229;
#20;
$display("Result = %d", result); assert(result ==556324);
row = 230;
#20;
$display("Result = %d", result); assert(result ==1820977);
row = 231;
#20;
$display("Result = %d", result); assert(result ==15286515);
row = 232;
#20;
$display("Result = %d", result); assert(result ==1028358);
row = 233;
#20;
$display("Result = %d", result); assert(result ==1543427);
row = 234;
#20;
$display("Result = %d", result); assert(result ==2192356);
row = 235;
#20;
$display("Result = %d", result); assert(result ==13652852);
row = 236;
#20;
$display("Result = %d", result); assert(result ==14069507);
row = 237;
#20;
$display("Result = %d", result); assert(result ==7573883);
row = 238;
#20;
$display("Result = %d", result); assert(result ==11701366);
row = 239;
#20;
$display("Result = %d", result); assert(result ==14610650);
row = 240;
#20;
$display("Result = %d", result); assert(result ==9578996);
row = 241;
#20;
$display("Result = %d", result); assert(result ==11623904);
row = 242;
#20;
$display("Result = %d", result); assert(result ==12429645);
row = 243;
#20;
$display("Result = %d", result); assert(result ==12492210);
row = 244;
#20;
$display("Result = %d", result); assert(result ==8301141);
row = 245;
#20;
$display("Result = %d", result); assert(result ==4607131);
row = 246;
#20;
$display("Result = %d", result); assert(result ==6180710);
row = 247;
#20;
$display("Result = %d", result); assert(result ==2022678);
row = 248;
#20;
$display("Result = %d", result); assert(result ==10821629);
row = 249;
#20;
$display("Result = %d", result); assert(result ==10451852);
row = 250;
#20;
$display("Result = %d", result); assert(result ==14112880);
row = 251;
#20;
$display("Result = %d", result); assert(result ==6090102);
row = 252;
#20;
$display("Result = %d", result); assert(result ==10848278);
row = 253;
#20;
$display("Result = %d", result); assert(result ==3543231);
row = 254;
#20;
$display("Result = %d", result); assert(result ==16590081);
row = 255;
#20;
$display("Result = %d", result); assert(result ==4044486);
row = 256;
#20;
$display("Result = %d", result); assert(result ==8698236);
en=0;
rst_n=0;
#100;
rst_n=1;
#100;
en=1;
#20;
ciphertext_select = 0;
row = 0;
ciphertext_entry =5642269;
#20;
row = 1;
ciphertext_entry =3086838;
#20;
row = 2;
ciphertext_entry =4398916;
#20;
row = 3;
ciphertext_entry =5056072;
#20;
row = 4;
ciphertext_entry =3101989;
#20;
row = 5;
ciphertext_entry =5323849;
#20;
row = 6;
ciphertext_entry =3017298;
#20;
row = 7;
ciphertext_entry =7869721;
#20;
row = 8;
ciphertext_entry =7148209;
#20;
row = 9;
ciphertext_entry =2237385;
#20;
row = 10;
ciphertext_entry =6619128;
#20;
row = 11;
ciphertext_entry =3379848;
#20;
row = 12;
ciphertext_entry =10488985;
#20;
row = 13;
ciphertext_entry =5364227;
#20;
row = 14;
ciphertext_entry =6797588;
#20;
row = 15;
ciphertext_entry =13625708;
#20;
row = 16;
ciphertext_entry =5471905;
#20;
row = 17;
ciphertext_entry =10692068;
#20;
row = 18;
ciphertext_entry =10000350;
#20;
row = 19;
ciphertext_entry =7096620;
#20;
row = 20;
ciphertext_entry =3181210;
#20;
row = 21;
ciphertext_entry =12223224;
#20;
row = 22;
ciphertext_entry =4867869;
#20;
row = 23;
ciphertext_entry =2646835;
#20;
row = 24;
ciphertext_entry =14545437;
#20;
row = 25;
ciphertext_entry =12887216;
#20;
row = 26;
ciphertext_entry =7428109;
#20;
row = 27;
ciphertext_entry =5922181;
#20;
row = 28;
ciphertext_entry =1226202;
#20;
row = 29;
ciphertext_entry =4757402;
#20;
row = 30;
ciphertext_entry =15576320;
#20;
row = 31;
ciphertext_entry =8242336;
#20;
row = 32;
ciphertext_entry =11104038;
#20;
row = 33;
ciphertext_entry =12648277;
#20;
row = 34;
ciphertext_entry =11512259;
#20;
row = 35;
ciphertext_entry =11861047;
#20;
row = 36;
ciphertext_entry =6827319;
#20;
row = 37;
ciphertext_entry =2855764;
#20;
row = 38;
ciphertext_entry =14355044;
#20;
row = 39;
ciphertext_entry =12255716;
#20;
row = 40;
ciphertext_entry =16421261;
#20;
row = 41;
ciphertext_entry =8530556;
#20;
row = 42;
ciphertext_entry =9088426;
#20;
row = 43;
ciphertext_entry =6880239;
#20;
row = 44;
ciphertext_entry =14401374;
#20;
row = 45;
ciphertext_entry =13905080;
#20;
row = 46;
ciphertext_entry =11418914;
#20;
row = 47;
ciphertext_entry =2719900;
#20;
row = 48;
ciphertext_entry =15448426;
#20;
row = 49;
ciphertext_entry =2864918;
#20;
row = 50;
ciphertext_entry =11383231;
#20;
row = 51;
ciphertext_entry =11415135;
#20;
row = 52;
ciphertext_entry =11555920;
#20;
row = 53;
ciphertext_entry =13716023;
#20;
row = 54;
ciphertext_entry =3957627;
#20;
row = 55;
ciphertext_entry =10312326;
#20;
row = 56;
ciphertext_entry =12174185;
#20;
row = 57;
ciphertext_entry =12073028;
#20;
row = 58;
ciphertext_entry =11876746;
#20;
row = 59;
ciphertext_entry =12786015;
#20;
row = 60;
ciphertext_entry =4814680;
#20;
row = 61;
ciphertext_entry =10525395;
#20;
row = 62;
ciphertext_entry =8349695;
#20;
row = 63;
ciphertext_entry =13984582;
#20;
row = 64;
ciphertext_entry =13057614;
#20;
row = 65;
ciphertext_entry =9652913;
#20;
row = 66;
ciphertext_entry =12061179;
#20;
row = 67;
ciphertext_entry =9115166;
#20;
row = 68;
ciphertext_entry =1045559;
#20;
row = 69;
ciphertext_entry =10581983;
#20;
row = 70;
ciphertext_entry =10673135;
#20;
row = 71;
ciphertext_entry =10908996;
#20;
row = 72;
ciphertext_entry =16007359;
#20;
row = 73;
ciphertext_entry =14660002;
#20;
row = 74;
ciphertext_entry =13979241;
#20;
row = 75;
ciphertext_entry =5380861;
#20;
row = 76;
ciphertext_entry =14292751;
#20;
row = 77;
ciphertext_entry =5358223;
#20;
row = 78;
ciphertext_entry =14865534;
#20;
row = 79;
ciphertext_entry =3261285;
#20;
row = 80;
ciphertext_entry =8820538;
#20;
row = 81;
ciphertext_entry =15406965;
#20;
row = 82;
ciphertext_entry =515576;
#20;
row = 83;
ciphertext_entry =15336274;
#20;
row = 84;
ciphertext_entry =4227748;
#20;
row = 85;
ciphertext_entry =10940536;
#20;
row = 86;
ciphertext_entry =15537510;
#20;
row = 87;
ciphertext_entry =15262270;
#20;
row = 88;
ciphertext_entry =16101356;
#20;
row = 89;
ciphertext_entry =4937333;
#20;
row = 90;
ciphertext_entry =12282975;
#20;
row = 91;
ciphertext_entry =5832144;
#20;
row = 92;
ciphertext_entry =4685901;
#20;
row = 93;
ciphertext_entry =13736852;
#20;
row = 94;
ciphertext_entry =14882910;
#20;
row = 95;
ciphertext_entry =11652248;
#20;
row = 96;
ciphertext_entry =5791352;
#20;
row = 97;
ciphertext_entry =10902292;
#20;
row = 98;
ciphertext_entry =10047326;
#20;
row = 99;
ciphertext_entry =2485678;
#20;
row = 100;
ciphertext_entry =5215655;
#20;
row = 101;
ciphertext_entry =1703647;
#20;
row = 102;
ciphertext_entry =11178922;
#20;
row = 103;
ciphertext_entry =2800619;
#20;
row = 104;
ciphertext_entry =13906880;
#20;
row = 105;
ciphertext_entry =12955023;
#20;
row = 106;
ciphertext_entry =858922;
#20;
row = 107;
ciphertext_entry =8491697;
#20;
row = 108;
ciphertext_entry =16089667;
#20;
row = 109;
ciphertext_entry =10004631;
#20;
row = 110;
ciphertext_entry =16480520;
#20;
row = 111;
ciphertext_entry =11183838;
#20;
row = 112;
ciphertext_entry =13152293;
#20;
row = 113;
ciphertext_entry =9189638;
#20;
row = 114;
ciphertext_entry =15818841;
#20;
row = 115;
ciphertext_entry =11025989;
#20;
row = 116;
ciphertext_entry =10220039;
#20;
row = 117;
ciphertext_entry =7136747;
#20;
row = 118;
ciphertext_entry =5569498;
#20;
row = 119;
ciphertext_entry =8053220;
#20;
row = 120;
ciphertext_entry =1070691;
#20;
row = 121;
ciphertext_entry =12464424;
#20;
row = 122;
ciphertext_entry =4888135;
#20;
row = 123;
ciphertext_entry =4352921;
#20;
row = 124;
ciphertext_entry =2727169;
#20;
row = 125;
ciphertext_entry =385162;
#20;
row = 126;
ciphertext_entry =10657542;
#20;
row = 127;
ciphertext_entry =12065756;
#20;
row = 128;
ciphertext_entry =164173;
#20;
ciphertext_select = 1;
row = 0;
ciphertext_entry =5642269;
#20;
$display("Result = %d", result); assert(result ==14663939);
row = 1;
ciphertext_entry =3086838;
#20;
$display("Result = %d", result); assert(result ==13952156);
row = 2;
ciphertext_entry =4398916;
#20;
$display("Result = %d", result); assert(result ==9927092);
row = 3;
ciphertext_entry =5056072;
#20;
$display("Result = %d", result); assert(result ==2104064);
row = 4;
ciphertext_entry =3101989;
#20;
$display("Result = %d", result); assert(result ==9085830);
row = 5;
ciphertext_entry =5323849;
#20;
$display("Result = %d", result); assert(result ==3394566);
row = 6;
ciphertext_entry =3017298;
#20;
$display("Result = %d", result); assert(result ==12694275);
row = 7;
ciphertext_entry =7869721;
#20;
$display("Result = %d", result); assert(result ==12014768);
row = 8;
ciphertext_entry =7148209;
#20;
$display("Result = %d", result); assert(result ==773870);
row = 9;
ciphertext_entry =2237385;
#20;
$display("Result = %d", result); assert(result ==6028400);
row = 10;
ciphertext_entry =6619128;
#20;
$display("Result = %d", result); assert(result ==1273698);
row = 11;
ciphertext_entry =3379848;
#20;
$display("Result = %d", result); assert(result ==3702041);
row = 12;
ciphertext_entry =10488985;
#20;
$display("Result = %d", result); assert(result ==2696093);
row = 13;
ciphertext_entry =5364227;
#20;
$display("Result = %d", result); assert(result ==14745831);
row = 14;
ciphertext_entry =6797588;
#20;
$display("Result = %d", result); assert(result ==12063668);
row = 15;
ciphertext_entry =13625708;
#20;
$display("Result = %d", result); assert(result ==3219000);
row = 16;
ciphertext_entry =5471905;
#20;
$display("Result = %d", result); assert(result ==11824189);
row = 17;
ciphertext_entry =10692068;
#20;
$display("Result = %d", result); assert(result ==9926357);
row = 18;
ciphertext_entry =10000350;
#20;
$display("Result = %d", result); assert(result ==799622);
row = 19;
ciphertext_entry =7096620;
#20;
$display("Result = %d", result); assert(result ==3188166);
row = 20;
ciphertext_entry =3181210;
#20;
$display("Result = %d", result); assert(result ==15307544);
row = 21;
ciphertext_entry =12223224;
#20;
$display("Result = %d", result); assert(result ==15691866);
row = 22;
ciphertext_entry =4867869;
#20;
$display("Result = %d", result); assert(result ==14684862);
row = 23;
ciphertext_entry =2646835;
#20;
$display("Result = %d", result); assert(result ==4546899);
row = 24;
ciphertext_entry =14545437;
#20;
$display("Result = %d", result); assert(result ==9406931);
row = 25;
ciphertext_entry =12887216;
#20;
$display("Result = %d", result); assert(result ==6922939);
row = 26;
ciphertext_entry =7428109;
#20;
$display("Result = %d", result); assert(result ==13828239);
row = 27;
ciphertext_entry =5922181;
#20;
$display("Result = %d", result); assert(result ==8729375);
row = 28;
ciphertext_entry =1226202;
#20;
$display("Result = %d", result); assert(result ==6209367);
row = 29;
ciphertext_entry =4757402;
#20;
$display("Result = %d", result); assert(result ==5424826);
row = 30;
ciphertext_entry =15576320;
#20;
$display("Result = %d", result); assert(result ==8958541);
row = 31;
ciphertext_entry =8242336;
#20;
$display("Result = %d", result); assert(result ==15329798);
row = 32;
ciphertext_entry =11104038;
#20;
$display("Result = %d", result); assert(result ==15306943);
row = 33;
ciphertext_entry =12648277;
#20;
$display("Result = %d", result); assert(result ==7592107);
row = 34;
ciphertext_entry =11512259;
#20;
$display("Result = %d", result); assert(result ==11056323);
row = 35;
ciphertext_entry =11861047;
#20;
$display("Result = %d", result); assert(result ==1446890);
row = 36;
ciphertext_entry =6827319;
#20;
$display("Result = %d", result); assert(result ==1113996);
row = 37;
ciphertext_entry =2855764;
#20;
$display("Result = %d", result); assert(result ==3429752);
row = 38;
ciphertext_entry =14355044;
#20;
$display("Result = %d", result); assert(result ==1639706);
row = 39;
ciphertext_entry =12255716;
#20;
$display("Result = %d", result); assert(result ==8545130);
row = 40;
ciphertext_entry =16421261;
#20;
$display("Result = %d", result); assert(result ==5078978);
row = 41;
ciphertext_entry =8530556;
#20;
$display("Result = %d", result); assert(result ==6574239);
row = 42;
ciphertext_entry =9088426;
#20;
$display("Result = %d", result); assert(result ==10681421);
row = 43;
ciphertext_entry =6880239;
#20;
$display("Result = %d", result); assert(result ==4699014);
row = 44;
ciphertext_entry =14401374;
#20;
$display("Result = %d", result); assert(result ==1752897);
row = 45;
ciphertext_entry =13905080;
#20;
$display("Result = %d", result); assert(result ==7727305);
row = 46;
ciphertext_entry =11418914;
#20;
$display("Result = %d", result); assert(result ==8024754);
row = 47;
ciphertext_entry =2719900;
#20;
$display("Result = %d", result); assert(result ==2967031);
row = 48;
ciphertext_entry =15448426;
#20;
$display("Result = %d", result); assert(result ==3845812);
row = 49;
ciphertext_entry =2864918;
#20;
$display("Result = %d", result); assert(result ==1927620);
row = 50;
ciphertext_entry =11383231;
#20;
$display("Result = %d", result); assert(result ==10769069);
row = 51;
ciphertext_entry =11415135;
#20;
$display("Result = %d", result); assert(result ==641470);
row = 52;
ciphertext_entry =11555920;
#20;
$display("Result = %d", result); assert(result ==12847349);
row = 53;
ciphertext_entry =13716023;
#20;
$display("Result = %d", result); assert(result ==5443403);
row = 54;
ciphertext_entry =3957627;
#20;
$display("Result = %d", result); assert(result ==14161717);
row = 55;
ciphertext_entry =10312326;
#20;
$display("Result = %d", result); assert(result ==7139659);
row = 56;
ciphertext_entry =12174185;
#20;
$display("Result = %d", result); assert(result ==13542520);
row = 57;
ciphertext_entry =12073028;
#20;
$display("Result = %d", result); assert(result ==6749965);
row = 58;
ciphertext_entry =11876746;
#20;
$display("Result = %d", result); assert(result ==15820721);
row = 59;
ciphertext_entry =12786015;
#20;
$display("Result = %d", result); assert(result ==8589441);
row = 60;
ciphertext_entry =4814680;
#20;
$display("Result = %d", result); assert(result ==2213600);
row = 61;
ciphertext_entry =10525395;
#20;
$display("Result = %d", result); assert(result ==14137482);
row = 62;
ciphertext_entry =8349695;
#20;
$display("Result = %d", result); assert(result ==3423672);
row = 63;
ciphertext_entry =13984582;
#20;
$display("Result = %d", result); assert(result ==1837170);
row = 64;
ciphertext_entry =13057614;
#20;
$display("Result = %d", result); assert(result ==15162791);
row = 65;
ciphertext_entry =9652913;
#20;
$display("Result = %d", result); assert(result ==11825062);
row = 66;
ciphertext_entry =12061179;
#20;
$display("Result = %d", result); assert(result ==16173937);
row = 67;
ciphertext_entry =9115166;
#20;
$display("Result = %d", result); assert(result ==9346583);
row = 68;
ciphertext_entry =1045559;
#20;
$display("Result = %d", result); assert(result ==12971427);
row = 69;
ciphertext_entry =10581983;
#20;
$display("Result = %d", result); assert(result ==1382657);
row = 70;
ciphertext_entry =10673135;
#20;
$display("Result = %d", result); assert(result ==3293203);
row = 71;
ciphertext_entry =10908996;
#20;
$display("Result = %d", result); assert(result ==9910401);
row = 72;
ciphertext_entry =16007359;
#20;
$display("Result = %d", result); assert(result ==8158411);
row = 73;
ciphertext_entry =14660002;
#20;
$display("Result = %d", result); assert(result ==9166577);
row = 74;
ciphertext_entry =13979241;
#20;
$display("Result = %d", result); assert(result ==3177207);
row = 75;
ciphertext_entry =5380861;
#20;
$display("Result = %d", result); assert(result ==6732170);
row = 76;
ciphertext_entry =14292751;
#20;
$display("Result = %d", result); assert(result ==6512601);
row = 77;
ciphertext_entry =5358223;
#20;
$display("Result = %d", result); assert(result ==4921568);
row = 78;
ciphertext_entry =14865534;
#20;
$display("Result = %d", result); assert(result ==4100901);
row = 79;
ciphertext_entry =3261285;
#20;
$display("Result = %d", result); assert(result ==1899952);
row = 80;
ciphertext_entry =8820538;
#20;
$display("Result = %d", result); assert(result ==5467310);
row = 81;
ciphertext_entry =15406965;
#20;
$display("Result = %d", result); assert(result ==13269032);
row = 82;
ciphertext_entry =515576;
#20;
$display("Result = %d", result); assert(result ==13896020);
row = 83;
ciphertext_entry =15336274;
#20;
$display("Result = %d", result); assert(result ==14326920);
row = 84;
ciphertext_entry =4227748;
#20;
$display("Result = %d", result); assert(result ==14502210);
row = 85;
ciphertext_entry =10940536;
#20;
$display("Result = %d", result); assert(result ==6304392);
row = 86;
ciphertext_entry =15537510;
#20;
$display("Result = %d", result); assert(result ==10634305);
row = 87;
ciphertext_entry =15262270;
#20;
$display("Result = %d", result); assert(result ==4979627);
row = 88;
ciphertext_entry =16101356;
#20;
$display("Result = %d", result); assert(result ==10462);
row = 89;
ciphertext_entry =4937333;
#20;
$display("Result = %d", result); assert(result ==8382718);
row = 90;
ciphertext_entry =12282975;
#20;
$display("Result = %d", result); assert(result ==13449115);
row = 91;
ciphertext_entry =5832144;
#20;
$display("Result = %d", result); assert(result ==13705307);
row = 92;
ciphertext_entry =4685901;
#20;
$display("Result = %d", result); assert(result ==2420486);
row = 93;
ciphertext_entry =13736852;
#20;
$display("Result = %d", result); assert(result ==15897284);
row = 94;
ciphertext_entry =14882910;
#20;
$display("Result = %d", result); assert(result ==9536294);
row = 95;
ciphertext_entry =11652248;
#20;
$display("Result = %d", result); assert(result ==15463837);
row = 96;
ciphertext_entry =5791352;
#20;
$display("Result = %d", result); assert(result ==6698986);
row = 97;
ciphertext_entry =10902292;
#20;
$display("Result = %d", result); assert(result ==448761);
row = 98;
ciphertext_entry =10047326;
#20;
$display("Result = %d", result); assert(result ==9255738);
row = 99;
ciphertext_entry =2485678;
#20;
$display("Result = %d", result); assert(result ==15176272);
row = 100;
ciphertext_entry =5215655;
#20;
$display("Result = %d", result); assert(result ==4271781);
row = 101;
ciphertext_entry =1703647;
#20;
$display("Result = %d", result); assert(result ==5354255);
row = 102;
ciphertext_entry =11178922;
#20;
$display("Result = %d", result); assert(result ==10556639);
row = 103;
ciphertext_entry =2800619;
#20;
$display("Result = %d", result); assert(result ==10057405);
row = 104;
ciphertext_entry =13906880;
#20;
$display("Result = %d", result); assert(result ==3610606);
row = 105;
ciphertext_entry =12955023;
#20;
$display("Result = %d", result); assert(result ==8028898);
row = 106;
ciphertext_entry =858922;
#20;
$display("Result = %d", result); assert(result ==13946955);
row = 107;
ciphertext_entry =8491697;
#20;
$display("Result = %d", result); assert(result ==9844852);
row = 108;
ciphertext_entry =16089667;
#20;
$display("Result = %d", result); assert(result ==3949826);
row = 109;
ciphertext_entry =10004631;
#20;
$display("Result = %d", result); assert(result ==16435605);
row = 110;
ciphertext_entry =16480520;
#20;
$display("Result = %d", result); assert(result ==6180254);
row = 111;
ciphertext_entry =11183838;
#20;
$display("Result = %d", result); assert(result ==10037353);
row = 112;
ciphertext_entry =13152293;
#20;
$display("Result = %d", result); assert(result ==16336314);
row = 113;
ciphertext_entry =9189638;
#20;
$display("Result = %d", result); assert(result ==10967391);
row = 114;
ciphertext_entry =15818841;
#20;
$display("Result = %d", result); assert(result ==13241510);
row = 115;
ciphertext_entry =11025989;
#20;
$display("Result = %d", result); assert(result ==11205497);
row = 116;
ciphertext_entry =10220039;
#20;
$display("Result = %d", result); assert(result ==11745390);
row = 117;
ciphertext_entry =7136747;
#20;
$display("Result = %d", result); assert(result ==11096401);
row = 118;
ciphertext_entry =5569498;
#20;
$display("Result = %d", result); assert(result ==4643569);
row = 119;
ciphertext_entry =8053220;
#20;
$display("Result = %d", result); assert(result ==2240304);
row = 120;
ciphertext_entry =1070691;
#20;
$display("Result = %d", result); assert(result ==14743989);
row = 121;
ciphertext_entry =12464424;
#20;
$display("Result = %d", result); assert(result ==3758356);
row = 122;
ciphertext_entry =4888135;
#20;
$display("Result = %d", result); assert(result ==10047764);
row = 123;
ciphertext_entry =4352921;
#20;
$display("Result = %d", result); assert(result ==11826019);
row = 124;
ciphertext_entry =2727169;
#20;
$display("Result = %d", result); assert(result ==2776380);
row = 125;
ciphertext_entry =385162;
#20;
$display("Result = %d", result); assert(result ==6988360);
row = 126;
ciphertext_entry =10657542;
#20;
$display("Result = %d", result); assert(result ==9140078);
row = 127;
ciphertext_entry =12065756;
#20;
$display("Result = %d", result); assert(result ==4487376);
row = 128;
ciphertext_entry =164173;
#20;
$display("Result = %d", result); assert(result ==7169268);
ciphertext_select = 0;
row = 129;
#20;
$display("Result = %d", result); assert(result ==5052296);
row = 130;
#20;
$display("Result = %d", result); assert(result ==11270021);
row = 131;
#20;
$display("Result = %d", result); assert(result ==12879228);
row = 132;
#20;
$display("Result = %d", result); assert(result ==9411225);
row = 133;
#20;
$display("Result = %d", result); assert(result ==13056492);
row = 134;
#20;
$display("Result = %d", result); assert(result ==3825524);
row = 135;
#20;
$display("Result = %d", result); assert(result ==7664373);
row = 136;
#20;
$display("Result = %d", result); assert(result ==388238);
row = 137;
#20;
$display("Result = %d", result); assert(result ==13874135);
row = 138;
#20;
$display("Result = %d", result); assert(result ==5673332);
row = 139;
#20;
$display("Result = %d", result); assert(result ==3164004);
row = 140;
#20;
$display("Result = %d", result); assert(result ==13274000);
row = 141;
#20;
$display("Result = %d", result); assert(result ==8196038);
row = 142;
#20;
$display("Result = %d", result); assert(result ==14429506);
row = 143;
#20;
$display("Result = %d", result); assert(result ==12971538);
row = 144;
#20;
$display("Result = %d", result); assert(result ==4520101);
row = 145;
#20;
$display("Result = %d", result); assert(result ==2890475);
row = 146;
#20;
$display("Result = %d", result); assert(result ==16402190);
row = 147;
#20;
$display("Result = %d", result); assert(result ==13541161);
row = 148;
#20;
$display("Result = %d", result); assert(result ==5190887);
row = 149;
#20;
$display("Result = %d", result); assert(result ==7930445);
row = 150;
#20;
$display("Result = %d", result); assert(result ==1151970);
row = 151;
#20;
$display("Result = %d", result); assert(result ==394940);
row = 152;
#20;
$display("Result = %d", result); assert(result ==3191108);
row = 153;
#20;
$display("Result = %d", result); assert(result ==10088470);
row = 154;
#20;
$display("Result = %d", result); assert(result ==13722300);
row = 155;
#20;
$display("Result = %d", result); assert(result ==10816944);
row = 156;
#20;
$display("Result = %d", result); assert(result ==7933907);
row = 157;
#20;
$display("Result = %d", result); assert(result ==2167565);
row = 158;
#20;
$display("Result = %d", result); assert(result ==7122547);
row = 159;
#20;
$display("Result = %d", result); assert(result ==6462149);
row = 160;
#20;
$display("Result = %d", result); assert(result ==16505043);
row = 161;
#20;
$display("Result = %d", result); assert(result ==4572172);
row = 162;
#20;
$display("Result = %d", result); assert(result ==15063988);
row = 163;
#20;
$display("Result = %d", result); assert(result ==10804531);
row = 164;
#20;
$display("Result = %d", result); assert(result ==11463681);
row = 165;
#20;
$display("Result = %d", result); assert(result ==231088);
row = 166;
#20;
$display("Result = %d", result); assert(result ==3518796);
row = 167;
#20;
$display("Result = %d", result); assert(result ==4780762);
row = 168;
#20;
$display("Result = %d", result); assert(result ==3255752);
row = 169;
#20;
$display("Result = %d", result); assert(result ==14961651);
row = 170;
#20;
$display("Result = %d", result); assert(result ==14545682);
row = 171;
#20;
$display("Result = %d", result); assert(result ==501215);
row = 172;
#20;
$display("Result = %d", result); assert(result ==1422523);
row = 173;
#20;
$display("Result = %d", result); assert(result ==11602211);
row = 174;
#20;
$display("Result = %d", result); assert(result ==10273744);
row = 175;
#20;
$display("Result = %d", result); assert(result ==10526859);
row = 176;
#20;
$display("Result = %d", result); assert(result ==10851345);
row = 177;
#20;
$display("Result = %d", result); assert(result ==10573789);
row = 178;
#20;
$display("Result = %d", result); assert(result ==1281554);
row = 179;
#20;
$display("Result = %d", result); assert(result ==15123937);
row = 180;
#20;
$display("Result = %d", result); assert(result ==6515791);
row = 181;
#20;
$display("Result = %d", result); assert(result ==3712576);
row = 182;
#20;
$display("Result = %d", result); assert(result ==5739919);
row = 183;
#20;
$display("Result = %d", result); assert(result ==16228712);
row = 184;
#20;
$display("Result = %d", result); assert(result ==1471307);
row = 185;
#20;
$display("Result = %d", result); assert(result ==8603342);
row = 186;
#20;
$display("Result = %d", result); assert(result ==14033414);
row = 187;
#20;
$display("Result = %d", result); assert(result ==2511213);
row = 188;
#20;
$display("Result = %d", result); assert(result ==14357821);
row = 189;
#20;
$display("Result = %d", result); assert(result ==15797272);
row = 190;
#20;
$display("Result = %d", result); assert(result ==14772726);
row = 191;
#20;
$display("Result = %d", result); assert(result ==15959437);
row = 192;
#20;
$display("Result = %d", result); assert(result ==2093983);
row = 193;
#20;
$display("Result = %d", result); assert(result ==10774010);
row = 194;
#20;
$display("Result = %d", result); assert(result ==11482724);
row = 195;
#20;
$display("Result = %d", result); assert(result ==2061331);
row = 196;
#20;
$display("Result = %d", result); assert(result ==10427655);
row = 197;
#20;
$display("Result = %d", result); assert(result ==1320450);
row = 198;
#20;
$display("Result = %d", result); assert(result ==6437525);
row = 199;
#20;
$display("Result = %d", result); assert(result ==3186622);
row = 200;
#20;
$display("Result = %d", result); assert(result ==3551081);
row = 201;
#20;
$display("Result = %d", result); assert(result ==15022238);
row = 202;
#20;
$display("Result = %d", result); assert(result ==5439264);
row = 203;
#20;
$display("Result = %d", result); assert(result ==1241020);
row = 204;
#20;
$display("Result = %d", result); assert(result ==3022910);
row = 205;
#20;
$display("Result = %d", result); assert(result ==9791610);
row = 206;
#20;
$display("Result = %d", result); assert(result ==6403304);
row = 207;
#20;
$display("Result = %d", result); assert(result ==14038202);
row = 208;
#20;
$display("Result = %d", result); assert(result ==13161080);
row = 209;
#20;
$display("Result = %d", result); assert(result ==2459445);
row = 210;
#20;
$display("Result = %d", result); assert(result ==803601);
row = 211;
#20;
$display("Result = %d", result); assert(result ==14231920);
row = 212;
#20;
$display("Result = %d", result); assert(result ==8101020);
row = 213;
#20;
$display("Result = %d", result); assert(result ==2339394);
row = 214;
#20;
$display("Result = %d", result); assert(result ==13647563);
row = 215;
#20;
$display("Result = %d", result); assert(result ==9885567);
row = 216;
#20;
$display("Result = %d", result); assert(result ==11342280);
row = 217;
#20;
$display("Result = %d", result); assert(result ==1204906);
row = 218;
#20;
$display("Result = %d", result); assert(result ==1052755);
row = 219;
#20;
$display("Result = %d", result); assert(result ==15809912);
row = 220;
#20;
$display("Result = %d", result); assert(result ==13996040);
row = 221;
#20;
$display("Result = %d", result); assert(result ==8866338);
row = 222;
#20;
$display("Result = %d", result); assert(result ==6578422);
row = 223;
#20;
$display("Result = %d", result); assert(result ==15274582);
row = 224;
#20;
$display("Result = %d", result); assert(result ==9393326);
row = 225;
#20;
$display("Result = %d", result); assert(result ==2988448);
row = 226;
#20;
$display("Result = %d", result); assert(result ==16311919);
row = 227;
#20;
$display("Result = %d", result); assert(result ==2012885);
row = 228;
#20;
$display("Result = %d", result); assert(result ==7962584);
row = 229;
#20;
$display("Result = %d", result); assert(result ==8107229);
row = 230;
#20;
$display("Result = %d", result); assert(result ==10670781);
row = 231;
#20;
$display("Result = %d", result); assert(result ==2792076);
row = 232;
#20;
$display("Result = %d", result); assert(result ==11277396);
row = 233;
#20;
$display("Result = %d", result); assert(result ==6337229);
row = 234;
#20;
$display("Result = %d", result); assert(result ==8508118);
row = 235;
#20;
$display("Result = %d", result); assert(result ==10887457);
row = 236;
#20;
$display("Result = %d", result); assert(result ==6702034);
row = 237;
#20;
$display("Result = %d", result); assert(result ==3873375);
row = 238;
#20;
$display("Result = %d", result); assert(result ==16438850);
row = 239;
#20;
$display("Result = %d", result); assert(result ==6755251);
row = 240;
#20;
$display("Result = %d", result); assert(result ==810250);
row = 241;
#20;
$display("Result = %d", result); assert(result ==6218645);
row = 242;
#20;
$display("Result = %d", result); assert(result ==10241);
row = 243;
#20;
$display("Result = %d", result); assert(result ==14817877);
row = 244;
#20;
$display("Result = %d", result); assert(result ==10908708);
row = 245;
#20;
$display("Result = %d", result); assert(result ==9173678);
row = 246;
#20;
$display("Result = %d", result); assert(result ==16418928);
row = 247;
#20;
$display("Result = %d", result); assert(result ==4157811);
row = 248;
#20;
$display("Result = %d", result); assert(result ==2939444);
row = 249;
#20;
$display("Result = %d", result); assert(result ==9985445);
row = 250;
#20;
$display("Result = %d", result); assert(result ==7961785);
row = 251;
#20;
$display("Result = %d", result); assert(result ==9713981);
row = 252;
#20;
$display("Result = %d", result); assert(result ==12253066);
row = 253;
#20;
$display("Result = %d", result); assert(result ==6145141);
row = 254;
#20;
$display("Result = %d", result); assert(result ==12886018);
row = 255;
#20;
$display("Result = %d", result); assert(result ==3819708);
row = 256;
#20;
$display("Result = %d", result); assert(result ==12392963);
en=0;
rst_n=0;
#100;
rst_n=1;
#100;
en=1;
#20;
ciphertext_select = 0;
row = 0;
ciphertext_entry =9183290;
#20;
row = 1;
ciphertext_entry =11535033;
#20;
row = 2;
ciphertext_entry =372367;
#20;
row = 3;
ciphertext_entry =12542413;
#20;
row = 4;
ciphertext_entry =7014866;
#20;
row = 5;
ciphertext_entry =8478507;
#20;
row = 6;
ciphertext_entry =8104661;
#20;
row = 7;
ciphertext_entry =7946179;
#20;
row = 8;
ciphertext_entry =5425860;
#20;
row = 9;
ciphertext_entry =8541055;
#20;
row = 10;
ciphertext_entry =15425745;
#20;
row = 11;
ciphertext_entry =16741112;
#20;
row = 12;
ciphertext_entry =3294334;
#20;
row = 13;
ciphertext_entry =2771410;
#20;
row = 14;
ciphertext_entry =12161558;
#20;
row = 15;
ciphertext_entry =1177176;
#20;
row = 16;
ciphertext_entry =11204810;
#20;
row = 17;
ciphertext_entry =13741981;
#20;
row = 18;
ciphertext_entry =8149671;
#20;
row = 19;
ciphertext_entry =9183388;
#20;
row = 20;
ciphertext_entry =14751153;
#20;
row = 21;
ciphertext_entry =698178;
#20;
row = 22;
ciphertext_entry =7932043;
#20;
row = 23;
ciphertext_entry =5705532;
#20;
row = 24;
ciphertext_entry =12890545;
#20;
row = 25;
ciphertext_entry =10618758;
#20;
row = 26;
ciphertext_entry =8913462;
#20;
row = 27;
ciphertext_entry =8564383;
#20;
row = 28;
ciphertext_entry =16174185;
#20;
row = 29;
ciphertext_entry =1412210;
#20;
row = 30;
ciphertext_entry =508436;
#20;
row = 31;
ciphertext_entry =9005972;
#20;
row = 32;
ciphertext_entry =7364722;
#20;
row = 33;
ciphertext_entry =1323555;
#20;
row = 34;
ciphertext_entry =6116676;
#20;
row = 35;
ciphertext_entry =8346415;
#20;
row = 36;
ciphertext_entry =14927864;
#20;
row = 37;
ciphertext_entry =1473447;
#20;
row = 38;
ciphertext_entry =939361;
#20;
row = 39;
ciphertext_entry =1988906;
#20;
row = 40;
ciphertext_entry =16727419;
#20;
row = 41;
ciphertext_entry =14980714;
#20;
row = 42;
ciphertext_entry =3822310;
#20;
row = 43;
ciphertext_entry =9290041;
#20;
row = 44;
ciphertext_entry =11725363;
#20;
row = 45;
ciphertext_entry =2619163;
#20;
row = 46;
ciphertext_entry =9511510;
#20;
row = 47;
ciphertext_entry =15696609;
#20;
row = 48;
ciphertext_entry =6665637;
#20;
row = 49;
ciphertext_entry =6353636;
#20;
row = 50;
ciphertext_entry =7051844;
#20;
row = 51;
ciphertext_entry =15902151;
#20;
row = 52;
ciphertext_entry =8420811;
#20;
row = 53;
ciphertext_entry =15766140;
#20;
row = 54;
ciphertext_entry =7298167;
#20;
row = 55;
ciphertext_entry =13182056;
#20;
row = 56;
ciphertext_entry =9327792;
#20;
row = 57;
ciphertext_entry =9303334;
#20;
row = 58;
ciphertext_entry =14379825;
#20;
row = 59;
ciphertext_entry =5613328;
#20;
row = 60;
ciphertext_entry =12979911;
#20;
row = 61;
ciphertext_entry =8103378;
#20;
row = 62;
ciphertext_entry =7351368;
#20;
row = 63;
ciphertext_entry =9003882;
#20;
row = 64;
ciphertext_entry =9393268;
#20;
row = 65;
ciphertext_entry =10409410;
#20;
row = 66;
ciphertext_entry =16167550;
#20;
row = 67;
ciphertext_entry =8065303;
#20;
row = 68;
ciphertext_entry =12449397;
#20;
row = 69;
ciphertext_entry =9782614;
#20;
row = 70;
ciphertext_entry =6768735;
#20;
row = 71;
ciphertext_entry =12496123;
#20;
row = 72;
ciphertext_entry =12443013;
#20;
row = 73;
ciphertext_entry =4330944;
#20;
row = 74;
ciphertext_entry =7996447;
#20;
row = 75;
ciphertext_entry =4690593;
#20;
row = 76;
ciphertext_entry =3921940;
#20;
row = 77;
ciphertext_entry =4528747;
#20;
row = 78;
ciphertext_entry =4424895;
#20;
row = 79;
ciphertext_entry =7672832;
#20;
row = 80;
ciphertext_entry =7305345;
#20;
row = 81;
ciphertext_entry =13883908;
#20;
row = 82;
ciphertext_entry =13728512;
#20;
row = 83;
ciphertext_entry =15360446;
#20;
row = 84;
ciphertext_entry =12644495;
#20;
row = 85;
ciphertext_entry =390060;
#20;
row = 86;
ciphertext_entry =5006431;
#20;
row = 87;
ciphertext_entry =2037621;
#20;
row = 88;
ciphertext_entry =7179676;
#20;
row = 89;
ciphertext_entry =1337286;
#20;
row = 90;
ciphertext_entry =12800410;
#20;
row = 91;
ciphertext_entry =2248403;
#20;
row = 92;
ciphertext_entry =10669948;
#20;
row = 93;
ciphertext_entry =8434134;
#20;
row = 94;
ciphertext_entry =1527198;
#20;
row = 95;
ciphertext_entry =12305619;
#20;
row = 96;
ciphertext_entry =16035573;
#20;
row = 97;
ciphertext_entry =4551789;
#20;
row = 98;
ciphertext_entry =15426971;
#20;
row = 99;
ciphertext_entry =10173033;
#20;
row = 100;
ciphertext_entry =527931;
#20;
row = 101;
ciphertext_entry =5734167;
#20;
row = 102;
ciphertext_entry =12404866;
#20;
row = 103;
ciphertext_entry =5473500;
#20;
row = 104;
ciphertext_entry =2997557;
#20;
row = 105;
ciphertext_entry =662520;
#20;
row = 106;
ciphertext_entry =14972561;
#20;
row = 107;
ciphertext_entry =7531406;
#20;
row = 108;
ciphertext_entry =13726406;
#20;
row = 109;
ciphertext_entry =7884913;
#20;
row = 110;
ciphertext_entry =8651350;
#20;
row = 111;
ciphertext_entry =2878371;
#20;
row = 112;
ciphertext_entry =6155427;
#20;
row = 113;
ciphertext_entry =2271846;
#20;
row = 114;
ciphertext_entry =3246871;
#20;
row = 115;
ciphertext_entry =805265;
#20;
row = 116;
ciphertext_entry =16471672;
#20;
row = 117;
ciphertext_entry =9295089;
#20;
row = 118;
ciphertext_entry =28867;
#20;
row = 119;
ciphertext_entry =6908596;
#20;
row = 120;
ciphertext_entry =3553164;
#20;
row = 121;
ciphertext_entry =6043564;
#20;
row = 122;
ciphertext_entry =7368226;
#20;
row = 123;
ciphertext_entry =15725853;
#20;
row = 124;
ciphertext_entry =3980842;
#20;
row = 125;
ciphertext_entry =1169678;
#20;
row = 126;
ciphertext_entry =16704076;
#20;
row = 127;
ciphertext_entry =6524549;
#20;
row = 128;
ciphertext_entry =15708200;
#20;
ciphertext_select = 1;
row = 0;
ciphertext_entry =9183290;
#20;
$display("Result = %d", result); assert(result ==13204434);
row = 1;
ciphertext_entry =11535033;
#20;
$display("Result = %d", result); assert(result ==10645223);
row = 2;
ciphertext_entry =372367;
#20;
$display("Result = %d", result); assert(result ==14342742);
row = 3;
ciphertext_entry =12542413;
#20;
$display("Result = %d", result); assert(result ==209605);
row = 4;
ciphertext_entry =7014866;
#20;
$display("Result = %d", result); assert(result ==7414751);
row = 5;
ciphertext_entry =8478507;
#20;
$display("Result = %d", result); assert(result ==954075);
row = 6;
ciphertext_entry =8104661;
#20;
$display("Result = %d", result); assert(result ==8068673);
row = 7;
ciphertext_entry =7946179;
#20;
$display("Result = %d", result); assert(result ==16446055);
row = 8;
ciphertext_entry =5425860;
#20;
$display("Result = %d", result); assert(result ==13881022);
row = 9;
ciphertext_entry =8541055;
#20;
$display("Result = %d", result); assert(result ==14667122);
row = 10;
ciphertext_entry =15425745;
#20;
$display("Result = %d", result); assert(result ==9290314);
row = 11;
ciphertext_entry =16741112;
#20;
$display("Result = %d", result); assert(result ==2077341);
row = 12;
ciphertext_entry =3294334;
#20;
$display("Result = %d", result); assert(result ==6569787);
row = 13;
ciphertext_entry =2771410;
#20;
$display("Result = %d", result); assert(result ==6573925);
row = 14;
ciphertext_entry =12161558;
#20;
$display("Result = %d", result); assert(result ==11014295);
row = 15;
ciphertext_entry =1177176;
#20;
$display("Result = %d", result); assert(result ==5989911);
row = 16;
ciphertext_entry =11204810;
#20;
$display("Result = %d", result); assert(result ==8947174);
row = 17;
ciphertext_entry =13741981;
#20;
$display("Result = %d", result); assert(result ==10415217);
row = 18;
ciphertext_entry =8149671;
#20;
$display("Result = %d", result); assert(result ==51254);
row = 19;
ciphertext_entry =9183388;
#20;
$display("Result = %d", result); assert(result ==14728793);
row = 20;
ciphertext_entry =14751153;
#20;
$display("Result = %d", result); assert(result ==12035341);
row = 21;
ciphertext_entry =698178;
#20;
$display("Result = %d", result); assert(result ==4653724);
row = 22;
ciphertext_entry =7932043;
#20;
$display("Result = %d", result); assert(result ==14391611);
row = 23;
ciphertext_entry =5705532;
#20;
$display("Result = %d", result); assert(result ==16301297);
row = 24;
ciphertext_entry =12890545;
#20;
$display("Result = %d", result); assert(result ==11328204);
row = 25;
ciphertext_entry =10618758;
#20;
$display("Result = %d", result); assert(result ==10908609);
row = 26;
ciphertext_entry =8913462;
#20;
$display("Result = %d", result); assert(result ==6462834);
row = 27;
ciphertext_entry =8564383;
#20;
$display("Result = %d", result); assert(result ==8533795);
row = 28;
ciphertext_entry =16174185;
#20;
$display("Result = %d", result); assert(result ==9978208);
row = 29;
ciphertext_entry =1412210;
#20;
$display("Result = %d", result); assert(result ==15923740);
row = 30;
ciphertext_entry =508436;
#20;
$display("Result = %d", result); assert(result ==1793012);
row = 31;
ciphertext_entry =9005972;
#20;
$display("Result = %d", result); assert(result ==13395202);
row = 32;
ciphertext_entry =7364722;
#20;
$display("Result = %d", result); assert(result ==4527924);
row = 33;
ciphertext_entry =1323555;
#20;
$display("Result = %d", result); assert(result ==8475669);
row = 34;
ciphertext_entry =6116676;
#20;
$display("Result = %d", result); assert(result ==5343612);
row = 35;
ciphertext_entry =8346415;
#20;
$display("Result = %d", result); assert(result ==15247676);
row = 36;
ciphertext_entry =14927864;
#20;
$display("Result = %d", result); assert(result ==2532257);
row = 37;
ciphertext_entry =1473447;
#20;
$display("Result = %d", result); assert(result ==16520944);
row = 38;
ciphertext_entry =939361;
#20;
$display("Result = %d", result); assert(result ==7917168);
row = 39;
ciphertext_entry =1988906;
#20;
$display("Result = %d", result); assert(result ==1983711);
row = 40;
ciphertext_entry =16727419;
#20;
$display("Result = %d", result); assert(result ==9068183);
row = 41;
ciphertext_entry =14980714;
#20;
$display("Result = %d", result); assert(result ==9267323);
row = 42;
ciphertext_entry =3822310;
#20;
$display("Result = %d", result); assert(result ==16404962);
row = 43;
ciphertext_entry =9290041;
#20;
$display("Result = %d", result); assert(result ==9378769);
row = 44;
ciphertext_entry =11725363;
#20;
$display("Result = %d", result); assert(result ==2527922);
row = 45;
ciphertext_entry =2619163;
#20;
$display("Result = %d", result); assert(result ==2099214);
row = 46;
ciphertext_entry =9511510;
#20;
$display("Result = %d", result); assert(result ==9366491);
row = 47;
ciphertext_entry =15696609;
#20;
$display("Result = %d", result); assert(result ==12635441);
row = 48;
ciphertext_entry =6665637;
#20;
$display("Result = %d", result); assert(result ==11900455);
row = 49;
ciphertext_entry =6353636;
#20;
$display("Result = %d", result); assert(result ==2922767);
row = 50;
ciphertext_entry =7051844;
#20;
$display("Result = %d", result); assert(result ==4629025);
row = 51;
ciphertext_entry =15902151;
#20;
$display("Result = %d", result); assert(result ==3898147);
row = 52;
ciphertext_entry =8420811;
#20;
$display("Result = %d", result); assert(result ==3159744);
row = 53;
ciphertext_entry =15766140;
#20;
$display("Result = %d", result); assert(result ==12980403);
row = 54;
ciphertext_entry =7298167;
#20;
$display("Result = %d", result); assert(result ==817177);
row = 55;
ciphertext_entry =13182056;
#20;
$display("Result = %d", result); assert(result ==9357258);
row = 56;
ciphertext_entry =9327792;
#20;
$display("Result = %d", result); assert(result ==15757208);
row = 57;
ciphertext_entry =9303334;
#20;
$display("Result = %d", result); assert(result ==8920651);
row = 58;
ciphertext_entry =14379825;
#20;
$display("Result = %d", result); assert(result ==6124283);
row = 59;
ciphertext_entry =5613328;
#20;
$display("Result = %d", result); assert(result ==8950237);
row = 60;
ciphertext_entry =12979911;
#20;
$display("Result = %d", result); assert(result ==113412);
row = 61;
ciphertext_entry =8103378;
#20;
$display("Result = %d", result); assert(result ==9106525);
row = 62;
ciphertext_entry =7351368;
#20;
$display("Result = %d", result); assert(result ==9868822);
row = 63;
ciphertext_entry =9003882;
#20;
$display("Result = %d", result); assert(result ==9070616);
row = 64;
ciphertext_entry =9393268;
#20;
$display("Result = %d", result); assert(result ==676770);
row = 65;
ciphertext_entry =10409410;
#20;
$display("Result = %d", result); assert(result ==14395627);
row = 66;
ciphertext_entry =16167550;
#20;
$display("Result = %d", result); assert(result ==560258);
row = 67;
ciphertext_entry =8065303;
#20;
$display("Result = %d", result); assert(result ==10457384);
row = 68;
ciphertext_entry =12449397;
#20;
$display("Result = %d", result); assert(result ==8182195);
row = 69;
ciphertext_entry =9782614;
#20;
$display("Result = %d", result); assert(result ==2338865);
row = 70;
ciphertext_entry =6768735;
#20;
$display("Result = %d", result); assert(result ==6940343);
row = 71;
ciphertext_entry =12496123;
#20;
$display("Result = %d", result); assert(result ==5574994);
row = 72;
ciphertext_entry =12443013;
#20;
$display("Result = %d", result); assert(result ==16056771);
row = 73;
ciphertext_entry =4330944;
#20;
$display("Result = %d", result); assert(result ==13665982);
row = 74;
ciphertext_entry =7996447;
#20;
$display("Result = %d", result); assert(result ==835197);
row = 75;
ciphertext_entry =4690593;
#20;
$display("Result = %d", result); assert(result ==16682778);
row = 76;
ciphertext_entry =3921940;
#20;
$display("Result = %d", result); assert(result ==2550864);
row = 77;
ciphertext_entry =4528747;
#20;
$display("Result = %d", result); assert(result ==16380271);
row = 78;
ciphertext_entry =4424895;
#20;
$display("Result = %d", result); assert(result ==9455643);
row = 79;
ciphertext_entry =7672832;
#20;
$display("Result = %d", result); assert(result ==10588106);
row = 80;
ciphertext_entry =7305345;
#20;
$display("Result = %d", result); assert(result ==2999103);
row = 81;
ciphertext_entry =13883908;
#20;
$display("Result = %d", result); assert(result ==7780941);
row = 82;
ciphertext_entry =13728512;
#20;
$display("Result = %d", result); assert(result ==1047474);
row = 83;
ciphertext_entry =15360446;
#20;
$display("Result = %d", result); assert(result ==2785021);
row = 84;
ciphertext_entry =12644495;
#20;
$display("Result = %d", result); assert(result ==12789644);
row = 85;
ciphertext_entry =390060;
#20;
$display("Result = %d", result); assert(result ==15775785);
row = 86;
ciphertext_entry =5006431;
#20;
$display("Result = %d", result); assert(result ==174639);
row = 87;
ciphertext_entry =2037621;
#20;
$display("Result = %d", result); assert(result ==4090398);
row = 88;
ciphertext_entry =7179676;
#20;
$display("Result = %d", result); assert(result ==13355675);
row = 89;
ciphertext_entry =1337286;
#20;
$display("Result = %d", result); assert(result ==12343392);
row = 90;
ciphertext_entry =12800410;
#20;
$display("Result = %d", result); assert(result ==10168489);
row = 91;
ciphertext_entry =2248403;
#20;
$display("Result = %d", result); assert(result ==5923477);
row = 92;
ciphertext_entry =10669948;
#20;
$display("Result = %d", result); assert(result ==14565492);
row = 93;
ciphertext_entry =8434134;
#20;
$display("Result = %d", result); assert(result ==13678878);
row = 94;
ciphertext_entry =1527198;
#20;
$display("Result = %d", result); assert(result ==16611846);
row = 95;
ciphertext_entry =12305619;
#20;
$display("Result = %d", result); assert(result ==9605442);
row = 96;
ciphertext_entry =16035573;
#20;
$display("Result = %d", result); assert(result ==10981162);
row = 97;
ciphertext_entry =4551789;
#20;
$display("Result = %d", result); assert(result ==8294805);
row = 98;
ciphertext_entry =15426971;
#20;
$display("Result = %d", result); assert(result ==11539719);
row = 99;
ciphertext_entry =10173033;
#20;
$display("Result = %d", result); assert(result ==11184042);
row = 100;
ciphertext_entry =527931;
#20;
$display("Result = %d", result); assert(result ==1354257);
row = 101;
ciphertext_entry =5734167;
#20;
$display("Result = %d", result); assert(result ==13463396);
row = 102;
ciphertext_entry =12404866;
#20;
$display("Result = %d", result); assert(result ==1133492);
row = 103;
ciphertext_entry =5473500;
#20;
$display("Result = %d", result); assert(result ==1533568);
row = 104;
ciphertext_entry =2997557;
#20;
$display("Result = %d", result); assert(result ==7484657);
row = 105;
ciphertext_entry =662520;
#20;
$display("Result = %d", result); assert(result ==8307894);
row = 106;
ciphertext_entry =14972561;
#20;
$display("Result = %d", result); assert(result ==15272834);
row = 107;
ciphertext_entry =7531406;
#20;
$display("Result = %d", result); assert(result ==1349829);
row = 108;
ciphertext_entry =13726406;
#20;
$display("Result = %d", result); assert(result ==1126629);
row = 109;
ciphertext_entry =7884913;
#20;
$display("Result = %d", result); assert(result ==3786784);
row = 110;
ciphertext_entry =8651350;
#20;
$display("Result = %d", result); assert(result ==11831960);
row = 111;
ciphertext_entry =2878371;
#20;
$display("Result = %d", result); assert(result ==4100898);
row = 112;
ciphertext_entry =6155427;
#20;
$display("Result = %d", result); assert(result ==690512);
row = 113;
ciphertext_entry =2271846;
#20;
$display("Result = %d", result); assert(result ==12573896);
row = 114;
ciphertext_entry =3246871;
#20;
$display("Result = %d", result); assert(result ==4129623);
row = 115;
ciphertext_entry =805265;
#20;
$display("Result = %d", result); assert(result ==13138224);
row = 116;
ciphertext_entry =16471672;
#20;
$display("Result = %d", result); assert(result ==14581642);
row = 117;
ciphertext_entry =9295089;
#20;
$display("Result = %d", result); assert(result ==12988744);
row = 118;
ciphertext_entry =28867;
#20;
$display("Result = %d", result); assert(result ==14237477);
row = 119;
ciphertext_entry =6908596;
#20;
$display("Result = %d", result); assert(result ==12863255);
row = 120;
ciphertext_entry =3553164;
#20;
$display("Result = %d", result); assert(result ==10736246);
row = 121;
ciphertext_entry =6043564;
#20;
$display("Result = %d", result); assert(result ==9372166);
row = 122;
ciphertext_entry =7368226;
#20;
$display("Result = %d", result); assert(result ==1374518);
row = 123;
ciphertext_entry =15725853;
#20;
$display("Result = %d", result); assert(result ==7274858);
row = 124;
ciphertext_entry =3980842;
#20;
$display("Result = %d", result); assert(result ==15076374);
row = 125;
ciphertext_entry =1169678;
#20;
$display("Result = %d", result); assert(result ==4109505);
row = 126;
ciphertext_entry =16704076;
#20;
$display("Result = %d", result); assert(result ==14630793);
row = 127;
ciphertext_entry =6524549;
#20;
$display("Result = %d", result); assert(result ==7258466);
row = 128;
ciphertext_entry =15708200;
#20;
$display("Result = %d", result); assert(result ==5076333);
ciphertext_select = 0;
row = 129;
#20;
$display("Result = %d", result); assert(result ==14950814);
row = 130;
#20;
$display("Result = %d", result); assert(result ==4167048);
row = 131;
#20;
$display("Result = %d", result); assert(result ==4073725);
row = 132;
#20;
$display("Result = %d", result); assert(result ==1333897);
row = 133;
#20;
$display("Result = %d", result); assert(result ==11593511);
row = 134;
#20;
$display("Result = %d", result); assert(result ==320907);
row = 135;
#20;
$display("Result = %d", result); assert(result ==1791752);
row = 136;
#20;
$display("Result = %d", result); assert(result ==3226440);
row = 137;
#20;
$display("Result = %d", result); assert(result ==12046756);
row = 138;
#20;
$display("Result = %d", result); assert(result ==8570110);
row = 139;
#20;
$display("Result = %d", result); assert(result ==5352181);
row = 140;
#20;
$display("Result = %d", result); assert(result ==15233552);
row = 141;
#20;
$display("Result = %d", result); assert(result ==11402992);
row = 142;
#20;
$display("Result = %d", result); assert(result ==3367103);
row = 143;
#20;
$display("Result = %d", result); assert(result ==5351);
row = 144;
#20;
$display("Result = %d", result); assert(result ==9613109);
row = 145;
#20;
$display("Result = %d", result); assert(result ==9871344);
row = 146;
#20;
$display("Result = %d", result); assert(result ==3296315);
row = 147;
#20;
$display("Result = %d", result); assert(result ==15050829);
row = 148;
#20;
$display("Result = %d", result); assert(result ==14585142);
row = 149;
#20;
$display("Result = %d", result); assert(result ==11471745);
row = 150;
#20;
$display("Result = %d", result); assert(result ==15503692);
row = 151;
#20;
$display("Result = %d", result); assert(result ==5437967);
row = 152;
#20;
$display("Result = %d", result); assert(result ==10112933);
row = 153;
#20;
$display("Result = %d", result); assert(result ==13190950);
row = 154;
#20;
$display("Result = %d", result); assert(result ==15391969);
row = 155;
#20;
$display("Result = %d", result); assert(result ==13040023);
row = 156;
#20;
$display("Result = %d", result); assert(result ==6701115);
row = 157;
#20;
$display("Result = %d", result); assert(result ==13891957);
row = 158;
#20;
$display("Result = %d", result); assert(result ==12038014);
row = 159;
#20;
$display("Result = %d", result); assert(result ==4466964);
row = 160;
#20;
$display("Result = %d", result); assert(result ==5276203);
row = 161;
#20;
$display("Result = %d", result); assert(result ==14673123);
row = 162;
#20;
$display("Result = %d", result); assert(result ==12084465);
row = 163;
#20;
$display("Result = %d", result); assert(result ==9906892);
row = 164;
#20;
$display("Result = %d", result); assert(result ==11415751);
row = 165;
#20;
$display("Result = %d", result); assert(result ==7577692);
row = 166;
#20;
$display("Result = %d", result); assert(result ==5821464);
row = 167;
#20;
$display("Result = %d", result); assert(result ==13002585);
row = 168;
#20;
$display("Result = %d", result); assert(result ==6270280);
row = 169;
#20;
$display("Result = %d", result); assert(result ==1657603);
row = 170;
#20;
$display("Result = %d", result); assert(result ==14319418);
row = 171;
#20;
$display("Result = %d", result); assert(result ==11231909);
row = 172;
#20;
$display("Result = %d", result); assert(result ==9081095);
row = 173;
#20;
$display("Result = %d", result); assert(result ==4592965);
row = 174;
#20;
$display("Result = %d", result); assert(result ==9850556);
row = 175;
#20;
$display("Result = %d", result); assert(result ==9047258);
row = 176;
#20;
$display("Result = %d", result); assert(result ==5700560);
row = 177;
#20;
$display("Result = %d", result); assert(result ==13783703);
row = 178;
#20;
$display("Result = %d", result); assert(result ==1575124);
row = 179;
#20;
$display("Result = %d", result); assert(result ==11220581);
row = 180;
#20;
$display("Result = %d", result); assert(result ==14605030);
row = 181;
#20;
$display("Result = %d", result); assert(result ==16572953);
row = 182;
#20;
$display("Result = %d", result); assert(result ==4479594);
row = 183;
#20;
$display("Result = %d", result); assert(result ==9669377);
row = 184;
#20;
$display("Result = %d", result); assert(result ==6238198);
row = 185;
#20;
$display("Result = %d", result); assert(result ==4983604);
row = 186;
#20;
$display("Result = %d", result); assert(result ==12321839);
row = 187;
#20;
$display("Result = %d", result); assert(result ==16400896);
row = 188;
#20;
$display("Result = %d", result); assert(result ==4147707);
row = 189;
#20;
$display("Result = %d", result); assert(result ==8700312);
row = 190;
#20;
$display("Result = %d", result); assert(result ==14893138);
row = 191;
#20;
$display("Result = %d", result); assert(result ==7287014);
row = 192;
#20;
$display("Result = %d", result); assert(result ==9551392);
row = 193;
#20;
$display("Result = %d", result); assert(result ==13951233);
row = 194;
#20;
$display("Result = %d", result); assert(result ==4128063);
row = 195;
#20;
$display("Result = %d", result); assert(result ==3125361);
row = 196;
#20;
$display("Result = %d", result); assert(result ==11979760);
row = 197;
#20;
$display("Result = %d", result); assert(result ==10614796);
row = 198;
#20;
$display("Result = %d", result); assert(result ==9017229);
row = 199;
#20;
$display("Result = %d", result); assert(result ==16667539);
row = 200;
#20;
$display("Result = %d", result); assert(result ==9356957);
row = 201;
#20;
$display("Result = %d", result); assert(result ==10683774);
row = 202;
#20;
$display("Result = %d", result); assert(result ==9136452);
row = 203;
#20;
$display("Result = %d", result); assert(result ==281050);
row = 204;
#20;
$display("Result = %d", result); assert(result ==6614043);
row = 205;
#20;
$display("Result = %d", result); assert(result ==7740925);
row = 206;
#20;
$display("Result = %d", result); assert(result ==10706697);
row = 207;
#20;
$display("Result = %d", result); assert(result ==5352264);
row = 208;
#20;
$display("Result = %d", result); assert(result ==369701);
row = 209;
#20;
$display("Result = %d", result); assert(result ==3234176);
row = 210;
#20;
$display("Result = %d", result); assert(result ==13381653);
row = 211;
#20;
$display("Result = %d", result); assert(result ==15906420);
row = 212;
#20;
$display("Result = %d", result); assert(result ==8296897);
row = 213;
#20;
$display("Result = %d", result); assert(result ==11888922);
row = 214;
#20;
$display("Result = %d", result); assert(result ==4189317);
row = 215;
#20;
$display("Result = %d", result); assert(result ==2924194);
row = 216;
#20;
$display("Result = %d", result); assert(result ==15396241);
row = 217;
#20;
$display("Result = %d", result); assert(result ==6714583);
row = 218;
#20;
$display("Result = %d", result); assert(result ==10103191);
row = 219;
#20;
$display("Result = %d", result); assert(result ==15694909);
row = 220;
#20;
$display("Result = %d", result); assert(result ==14828632);
row = 221;
#20;
$display("Result = %d", result); assert(result ==11344084);
row = 222;
#20;
$display("Result = %d", result); assert(result ==4802847);
row = 223;
#20;
$display("Result = %d", result); assert(result ==3210794);
row = 224;
#20;
$display("Result = %d", result); assert(result ==1329091);
row = 225;
#20;
$display("Result = %d", result); assert(result ==7690731);
row = 226;
#20;
$display("Result = %d", result); assert(result ==4169298);
row = 227;
#20;
$display("Result = %d", result); assert(result ==11455573);
row = 228;
#20;
$display("Result = %d", result); assert(result ==7983915);
row = 229;
#20;
$display("Result = %d", result); assert(result ==4355577);
row = 230;
#20;
$display("Result = %d", result); assert(result ==5885180);
row = 231;
#20;
$display("Result = %d", result); assert(result ==3676000);
row = 232;
#20;
$display("Result = %d", result); assert(result ==587728);
row = 233;
#20;
$display("Result = %d", result); assert(result ==2379874);
row = 234;
#20;
$display("Result = %d", result); assert(result ==6347403);
row = 235;
#20;
$display("Result = %d", result); assert(result ==14663201);
row = 236;
#20;
$display("Result = %d", result); assert(result ==7595459);
row = 237;
#20;
$display("Result = %d", result); assert(result ==10580230);
row = 238;
#20;
$display("Result = %d", result); assert(result ==16608558);
row = 239;
#20;
$display("Result = %d", result); assert(result ==9815950);
row = 240;
#20;
$display("Result = %d", result); assert(result ==14579043);
row = 241;
#20;
$display("Result = %d", result); assert(result ==9186024);
row = 242;
#20;
$display("Result = %d", result); assert(result ==1584212);
row = 243;
#20;
$display("Result = %d", result); assert(result ==11282587);
row = 244;
#20;
$display("Result = %d", result); assert(result ==6909149);
row = 245;
#20;
$display("Result = %d", result); assert(result ==1247275);
row = 246;
#20;
$display("Result = %d", result); assert(result ==4437868);
row = 247;
#20;
$display("Result = %d", result); assert(result ==11414939);
row = 248;
#20;
$display("Result = %d", result); assert(result ==10037488);
row = 249;
#20;
$display("Result = %d", result); assert(result ==7174961);
row = 250;
#20;
$display("Result = %d", result); assert(result ==6456889);
row = 251;
#20;
$display("Result = %d", result); assert(result ==14714032);
row = 252;
#20;
$display("Result = %d", result); assert(result ==11360996);
row = 253;
#20;
$display("Result = %d", result); assert(result ==651025);
row = 254;
#20;
$display("Result = %d", result); assert(result ==8859565);
row = 255;
#20;
$display("Result = %d", result); assert(result ==3430163);
row = 256;
#20;
$display("Result = %d", result); assert(result ==8803416);
en=0;
rst_n=0;
#100;
rst_n=1;
#100;
en=1;
#20;
ciphertext_select = 0;
row = 0;
ciphertext_entry =4670736;
#20;
row = 1;
ciphertext_entry =8861663;
#20;
row = 2;
ciphertext_entry =13093436;
#20;
row = 3;
ciphertext_entry =14915754;
#20;
row = 4;
ciphertext_entry =885301;
#20;
row = 5;
ciphertext_entry =11813896;
#20;
row = 6;
ciphertext_entry =1966680;
#20;
row = 7;
ciphertext_entry =8285649;
#20;
row = 8;
ciphertext_entry =14564978;
#20;
row = 9;
ciphertext_entry =13677681;
#20;
row = 10;
ciphertext_entry =10391871;
#20;
row = 11;
ciphertext_entry =16257447;
#20;
row = 12;
ciphertext_entry =13749331;
#20;
row = 13;
ciphertext_entry =11204574;
#20;
row = 14;
ciphertext_entry =5622369;
#20;
row = 15;
ciphertext_entry =13590102;
#20;
row = 16;
ciphertext_entry =12472781;
#20;
row = 17;
ciphertext_entry =14268626;
#20;
row = 18;
ciphertext_entry =6125388;
#20;
row = 19;
ciphertext_entry =11856754;
#20;
row = 20;
ciphertext_entry =13715153;
#20;
row = 21;
ciphertext_entry =11264711;
#20;
row = 22;
ciphertext_entry =9034324;
#20;
row = 23;
ciphertext_entry =10051387;
#20;
row = 24;
ciphertext_entry =16187766;
#20;
row = 25;
ciphertext_entry =10124067;
#20;
row = 26;
ciphertext_entry =15507996;
#20;
row = 27;
ciphertext_entry =15303470;
#20;
row = 28;
ciphertext_entry =4608851;
#20;
row = 29;
ciphertext_entry =671611;
#20;
row = 30;
ciphertext_entry =13049661;
#20;
row = 31;
ciphertext_entry =8164116;
#20;
row = 32;
ciphertext_entry =11683536;
#20;
row = 33;
ciphertext_entry =8148938;
#20;
row = 34;
ciphertext_entry =16279164;
#20;
row = 35;
ciphertext_entry =11687494;
#20;
row = 36;
ciphertext_entry =4462393;
#20;
row = 37;
ciphertext_entry =5065974;
#20;
row = 38;
ciphertext_entry =10466793;
#20;
row = 39;
ciphertext_entry =1283054;
#20;
row = 40;
ciphertext_entry =3037337;
#20;
row = 41;
ciphertext_entry =777635;
#20;
row = 42;
ciphertext_entry =11808773;
#20;
row = 43;
ciphertext_entry =14974759;
#20;
row = 44;
ciphertext_entry =7261564;
#20;
row = 45;
ciphertext_entry =8229925;
#20;
row = 46;
ciphertext_entry =13526394;
#20;
row = 47;
ciphertext_entry =12460809;
#20;
row = 48;
ciphertext_entry =15052294;
#20;
row = 49;
ciphertext_entry =16685683;
#20;
row = 50;
ciphertext_entry =5028070;
#20;
row = 51;
ciphertext_entry =5922914;
#20;
row = 52;
ciphertext_entry =6297372;
#20;
row = 53;
ciphertext_entry =8695580;
#20;
row = 54;
ciphertext_entry =14108986;
#20;
row = 55;
ciphertext_entry =12931592;
#20;
row = 56;
ciphertext_entry =10659046;
#20;
row = 57;
ciphertext_entry =5771915;
#20;
row = 58;
ciphertext_entry =11117053;
#20;
row = 59;
ciphertext_entry =8971090;
#20;
row = 60;
ciphertext_entry =412381;
#20;
row = 61;
ciphertext_entry =15452044;
#20;
row = 62;
ciphertext_entry =3175565;
#20;
row = 63;
ciphertext_entry =94091;
#20;
row = 64;
ciphertext_entry =15715466;
#20;
row = 65;
ciphertext_entry =5063375;
#20;
row = 66;
ciphertext_entry =15244781;
#20;
row = 67;
ciphertext_entry =2141011;
#20;
row = 68;
ciphertext_entry =8158460;
#20;
row = 69;
ciphertext_entry =8354541;
#20;
row = 70;
ciphertext_entry =7945145;
#20;
row = 71;
ciphertext_entry =2451926;
#20;
row = 72;
ciphertext_entry =5492431;
#20;
row = 73;
ciphertext_entry =6270281;
#20;
row = 74;
ciphertext_entry =3374093;
#20;
row = 75;
ciphertext_entry =597819;
#20;
row = 76;
ciphertext_entry =9318833;
#20;
row = 77;
ciphertext_entry =16155775;
#20;
row = 78;
ciphertext_entry =7285469;
#20;
row = 79;
ciphertext_entry =7767504;
#20;
row = 80;
ciphertext_entry =8975752;
#20;
row = 81;
ciphertext_entry =15485818;
#20;
row = 82;
ciphertext_entry =3501553;
#20;
row = 83;
ciphertext_entry =4758484;
#20;
row = 84;
ciphertext_entry =6581426;
#20;
row = 85;
ciphertext_entry =9036514;
#20;
row = 86;
ciphertext_entry =12371712;
#20;
row = 87;
ciphertext_entry =7407448;
#20;
row = 88;
ciphertext_entry =12515029;
#20;
row = 89;
ciphertext_entry =7970250;
#20;
row = 90;
ciphertext_entry =10526160;
#20;
row = 91;
ciphertext_entry =6706932;
#20;
row = 92;
ciphertext_entry =15993295;
#20;
row = 93;
ciphertext_entry =2137088;
#20;
row = 94;
ciphertext_entry =467546;
#20;
row = 95;
ciphertext_entry =5605666;
#20;
row = 96;
ciphertext_entry =2850830;
#20;
row = 97;
ciphertext_entry =15595093;
#20;
row = 98;
ciphertext_entry =13138120;
#20;
row = 99;
ciphertext_entry =4554535;
#20;
row = 100;
ciphertext_entry =734256;
#20;
row = 101;
ciphertext_entry =5805692;
#20;
row = 102;
ciphertext_entry =5451957;
#20;
row = 103;
ciphertext_entry =13096827;
#20;
row = 104;
ciphertext_entry =4260172;
#20;
row = 105;
ciphertext_entry =13396514;
#20;
row = 106;
ciphertext_entry =16680876;
#20;
row = 107;
ciphertext_entry =6722048;
#20;
row = 108;
ciphertext_entry =2834274;
#20;
row = 109;
ciphertext_entry =14511046;
#20;
row = 110;
ciphertext_entry =15404940;
#20;
row = 111;
ciphertext_entry =15007265;
#20;
row = 112;
ciphertext_entry =12545968;
#20;
row = 113;
ciphertext_entry =2176121;
#20;
row = 114;
ciphertext_entry =10812240;
#20;
row = 115;
ciphertext_entry =14216943;
#20;
row = 116;
ciphertext_entry =14341961;
#20;
row = 117;
ciphertext_entry =3124841;
#20;
row = 118;
ciphertext_entry =3246222;
#20;
row = 119;
ciphertext_entry =6464138;
#20;
row = 120;
ciphertext_entry =13405847;
#20;
row = 121;
ciphertext_entry =13433205;
#20;
row = 122;
ciphertext_entry =8678602;
#20;
row = 123;
ciphertext_entry =15433985;
#20;
row = 124;
ciphertext_entry =5716110;
#20;
row = 125;
ciphertext_entry =157732;
#20;
row = 126;
ciphertext_entry =8883810;
#20;
row = 127;
ciphertext_entry =14103754;
#20;
row = 128;
ciphertext_entry =5606096;
#20;
ciphertext_select = 1;
row = 0;
ciphertext_entry =4670736;
#20;
$display("Result = %d", result); assert(result ==12672976);
row = 1;
ciphertext_entry =8861663;
#20;
$display("Result = %d", result); assert(result ==3757683);
row = 2;
ciphertext_entry =13093436;
#20;
$display("Result = %d", result); assert(result ==13085036);
row = 3;
ciphertext_entry =14915754;
#20;
$display("Result = %d", result); assert(result ==6683664);
row = 4;
ciphertext_entry =885301;
#20;
$display("Result = %d", result); assert(result ==12898457);
row = 5;
ciphertext_entry =11813896;
#20;
$display("Result = %d", result); assert(result ==16679233);
row = 6;
ciphertext_entry =1966680;
#20;
$display("Result = %d", result); assert(result ==9586631);
row = 7;
ciphertext_entry =8285649;
#20;
$display("Result = %d", result); assert(result ==13485156);
row = 8;
ciphertext_entry =14564978;
#20;
$display("Result = %d", result); assert(result ==2517772);
row = 9;
ciphertext_entry =13677681;
#20;
$display("Result = %d", result); assert(result ==15773875);
row = 10;
ciphertext_entry =10391871;
#20;
$display("Result = %d", result); assert(result ==9782518);
row = 11;
ciphertext_entry =16257447;
#20;
$display("Result = %d", result); assert(result ==12698515);
row = 12;
ciphertext_entry =13749331;
#20;
$display("Result = %d", result); assert(result ==4557158);
row = 13;
ciphertext_entry =11204574;
#20;
$display("Result = %d", result); assert(result ==10973894);
row = 14;
ciphertext_entry =5622369;
#20;
$display("Result = %d", result); assert(result ==2446125);
row = 15;
ciphertext_entry =13590102;
#20;
$display("Result = %d", result); assert(result ==7253425);
row = 16;
ciphertext_entry =12472781;
#20;
$display("Result = %d", result); assert(result ==7595132);
row = 17;
ciphertext_entry =14268626;
#20;
$display("Result = %d", result); assert(result ==4903608);
row = 18;
ciphertext_entry =6125388;
#20;
$display("Result = %d", result); assert(result ==605881);
row = 19;
ciphertext_entry =11856754;
#20;
$display("Result = %d", result); assert(result ==12930895);
row = 20;
ciphertext_entry =13715153;
#20;
$display("Result = %d", result); assert(result ==11369266);
row = 21;
ciphertext_entry =11264711;
#20;
$display("Result = %d", result); assert(result ==4834245);
row = 22;
ciphertext_entry =9034324;
#20;
$display("Result = %d", result); assert(result ==14799724);
row = 23;
ciphertext_entry =10051387;
#20;
$display("Result = %d", result); assert(result ==16628769);
row = 24;
ciphertext_entry =16187766;
#20;
$display("Result = %d", result); assert(result ==1285071);
row = 25;
ciphertext_entry =10124067;
#20;
$display("Result = %d", result); assert(result ==14425677);
row = 26;
ciphertext_entry =15507996;
#20;
$display("Result = %d", result); assert(result ==9571773);
row = 27;
ciphertext_entry =15303470;
#20;
$display("Result = %d", result); assert(result ==9421693);
row = 28;
ciphertext_entry =4608851;
#20;
$display("Result = %d", result); assert(result ==3660537);
row = 29;
ciphertext_entry =671611;
#20;
$display("Result = %d", result); assert(result ==2379162);
row = 30;
ciphertext_entry =13049661;
#20;
$display("Result = %d", result); assert(result ==6056081);
row = 31;
ciphertext_entry =8164116;
#20;
$display("Result = %d", result); assert(result ==5193183);
row = 32;
ciphertext_entry =11683536;
#20;
$display("Result = %d", result); assert(result ==4942194);
row = 33;
ciphertext_entry =8148938;
#20;
$display("Result = %d", result); assert(result ==11387150);
row = 34;
ciphertext_entry =16279164;
#20;
$display("Result = %d", result); assert(result ==1276465);
row = 35;
ciphertext_entry =11687494;
#20;
$display("Result = %d", result); assert(result ==13645028);
row = 36;
ciphertext_entry =4462393;
#20;
$display("Result = %d", result); assert(result ==2692321);
row = 37;
ciphertext_entry =5065974;
#20;
$display("Result = %d", result); assert(result ==6562869);
row = 38;
ciphertext_entry =10466793;
#20;
$display("Result = %d", result); assert(result ==9913033);
row = 39;
ciphertext_entry =1283054;
#20;
$display("Result = %d", result); assert(result ==3697264);
row = 40;
ciphertext_entry =3037337;
#20;
$display("Result = %d", result); assert(result ==14663141);
row = 41;
ciphertext_entry =777635;
#20;
$display("Result = %d", result); assert(result ==3106043);
row = 42;
ciphertext_entry =11808773;
#20;
$display("Result = %d", result); assert(result ==5945243);
row = 43;
ciphertext_entry =14974759;
#20;
$display("Result = %d", result); assert(result ==7034174);
row = 44;
ciphertext_entry =7261564;
#20;
$display("Result = %d", result); assert(result ==2208965);
row = 45;
ciphertext_entry =8229925;
#20;
$display("Result = %d", result); assert(result ==7840114);
row = 46;
ciphertext_entry =13526394;
#20;
$display("Result = %d", result); assert(result ==11536126);
row = 47;
ciphertext_entry =12460809;
#20;
$display("Result = %d", result); assert(result ==8284139);
row = 48;
ciphertext_entry =15052294;
#20;
$display("Result = %d", result); assert(result ==1376812);
row = 49;
ciphertext_entry =16685683;
#20;
$display("Result = %d", result); assert(result ==8624906);
row = 50;
ciphertext_entry =5028070;
#20;
$display("Result = %d", result); assert(result ==8836970);
row = 51;
ciphertext_entry =5922914;
#20;
$display("Result = %d", result); assert(result ==7995330);
row = 52;
ciphertext_entry =6297372;
#20;
$display("Result = %d", result); assert(result ==8828333);
row = 53;
ciphertext_entry =8695580;
#20;
$display("Result = %d", result); assert(result ==772117);
row = 54;
ciphertext_entry =14108986;
#20;
$display("Result = %d", result); assert(result ==467032);
row = 55;
ciphertext_entry =12931592;
#20;
$display("Result = %d", result); assert(result ==16682490);
row = 56;
ciphertext_entry =10659046;
#20;
$display("Result = %d", result); assert(result ==13634218);
row = 57;
ciphertext_entry =5771915;
#20;
$display("Result = %d", result); assert(result ==308215);
row = 58;
ciphertext_entry =11117053;
#20;
$display("Result = %d", result); assert(result ==7830888);
row = 59;
ciphertext_entry =8971090;
#20;
$display("Result = %d", result); assert(result ==14928877);
row = 60;
ciphertext_entry =412381;
#20;
$display("Result = %d", result); assert(result ==5213055);
row = 61;
ciphertext_entry =15452044;
#20;
$display("Result = %d", result); assert(result ==2395499);
row = 62;
ciphertext_entry =3175565;
#20;
$display("Result = %d", result); assert(result ==1015959);
row = 63;
ciphertext_entry =94091;
#20;
$display("Result = %d", result); assert(result ==8979588);
row = 64;
ciphertext_entry =15715466;
#20;
$display("Result = %d", result); assert(result ==10806917);
row = 65;
ciphertext_entry =5063375;
#20;
$display("Result = %d", result); assert(result ==8426356);
row = 66;
ciphertext_entry =15244781;
#20;
$display("Result = %d", result); assert(result ==7552730);
row = 67;
ciphertext_entry =2141011;
#20;
$display("Result = %d", result); assert(result ==11014618);
row = 68;
ciphertext_entry =8158460;
#20;
$display("Result = %d", result); assert(result ==5917780);
row = 69;
ciphertext_entry =8354541;
#20;
$display("Result = %d", result); assert(result ==13294248);
row = 70;
ciphertext_entry =7945145;
#20;
$display("Result = %d", result); assert(result ==10096191);
row = 71;
ciphertext_entry =2451926;
#20;
$display("Result = %d", result); assert(result ==10011465);
row = 72;
ciphertext_entry =5492431;
#20;
$display("Result = %d", result); assert(result ==14689697);
row = 73;
ciphertext_entry =6270281;
#20;
$display("Result = %d", result); assert(result ==12265022);
row = 74;
ciphertext_entry =3374093;
#20;
$display("Result = %d", result); assert(result ==3063600);
row = 75;
ciphertext_entry =597819;
#20;
$display("Result = %d", result); assert(result ==13746676);
row = 76;
ciphertext_entry =9318833;
#20;
$display("Result = %d", result); assert(result ==5984285);
row = 77;
ciphertext_entry =16155775;
#20;
$display("Result = %d", result); assert(result ==4978661);
row = 78;
ciphertext_entry =7285469;
#20;
$display("Result = %d", result); assert(result ==10696173);
row = 79;
ciphertext_entry =7767504;
#20;
$display("Result = %d", result); assert(result ==9337903);
row = 80;
ciphertext_entry =8975752;
#20;
$display("Result = %d", result); assert(result ==4103061);
row = 81;
ciphertext_entry =15485818;
#20;
$display("Result = %d", result); assert(result ==12760654);
row = 82;
ciphertext_entry =3501553;
#20;
$display("Result = %d", result); assert(result ==15332911);
row = 83;
ciphertext_entry =4758484;
#20;
$display("Result = %d", result); assert(result ==7467651);
row = 84;
ciphertext_entry =6581426;
#20;
$display("Result = %d", result); assert(result ==14665281);
row = 85;
ciphertext_entry =9036514;
#20;
$display("Result = %d", result); assert(result ==5333137);
row = 86;
ciphertext_entry =12371712;
#20;
$display("Result = %d", result); assert(result ==4312332);
row = 87;
ciphertext_entry =7407448;
#20;
$display("Result = %d", result); assert(result ==6581563);
row = 88;
ciphertext_entry =12515029;
#20;
$display("Result = %d", result); assert(result ==12261887);
row = 89;
ciphertext_entry =7970250;
#20;
$display("Result = %d", result); assert(result ==14617992);
row = 90;
ciphertext_entry =10526160;
#20;
$display("Result = %d", result); assert(result ==15045084);
row = 91;
ciphertext_entry =6706932;
#20;
$display("Result = %d", result); assert(result ==1304580);
row = 92;
ciphertext_entry =15993295;
#20;
$display("Result = %d", result); assert(result ==13990937);
row = 93;
ciphertext_entry =2137088;
#20;
$display("Result = %d", result); assert(result ==7675833);
row = 94;
ciphertext_entry =467546;
#20;
$display("Result = %d", result); assert(result ==6386988);
row = 95;
ciphertext_entry =5605666;
#20;
$display("Result = %d", result); assert(result ==13530595);
row = 96;
ciphertext_entry =2850830;
#20;
$display("Result = %d", result); assert(result ==7506885);
row = 97;
ciphertext_entry =15595093;
#20;
$display("Result = %d", result); assert(result ==10392136);
row = 98;
ciphertext_entry =13138120;
#20;
$display("Result = %d", result); assert(result ==15607080);
row = 99;
ciphertext_entry =4554535;
#20;
$display("Result = %d", result); assert(result ==11721138);
row = 100;
ciphertext_entry =734256;
#20;
$display("Result = %d", result); assert(result ==15798798);
row = 101;
ciphertext_entry =5805692;
#20;
$display("Result = %d", result); assert(result ==15744310);
row = 102;
ciphertext_entry =5451957;
#20;
$display("Result = %d", result); assert(result ==15361546);
row = 103;
ciphertext_entry =13096827;
#20;
$display("Result = %d", result); assert(result ==12101675);
row = 104;
ciphertext_entry =4260172;
#20;
$display("Result = %d", result); assert(result ==12311929);
row = 105;
ciphertext_entry =13396514;
#20;
$display("Result = %d", result); assert(result ==15286361);
row = 106;
ciphertext_entry =16680876;
#20;
$display("Result = %d", result); assert(result ==8131554);
row = 107;
ciphertext_entry =6722048;
#20;
$display("Result = %d", result); assert(result ==137552);
row = 108;
ciphertext_entry =2834274;
#20;
$display("Result = %d", result); assert(result ==2209837);
row = 109;
ciphertext_entry =14511046;
#20;
$display("Result = %d", result); assert(result ==12430557);
row = 110;
ciphertext_entry =15404940;
#20;
$display("Result = %d", result); assert(result ==5038150);
row = 111;
ciphertext_entry =15007265;
#20;
$display("Result = %d", result); assert(result ==5266260);
row = 112;
ciphertext_entry =12545968;
#20;
$display("Result = %d", result); assert(result ==15169897);
row = 113;
ciphertext_entry =2176121;
#20;
$display("Result = %d", result); assert(result ==16443161);
row = 114;
ciphertext_entry =10812240;
#20;
$display("Result = %d", result); assert(result ==100332);
row = 115;
ciphertext_entry =14216943;
#20;
$display("Result = %d", result); assert(result ==5059226);
row = 116;
ciphertext_entry =14341961;
#20;
$display("Result = %d", result); assert(result ==13693289);
row = 117;
ciphertext_entry =3124841;
#20;
$display("Result = %d", result); assert(result ==1782155);
row = 118;
ciphertext_entry =3246222;
#20;
$display("Result = %d", result); assert(result ==2090202);
row = 119;
ciphertext_entry =6464138;
#20;
$display("Result = %d", result); assert(result ==15710088);
row = 120;
ciphertext_entry =13405847;
#20;
$display("Result = %d", result); assert(result ==1776365);
row = 121;
ciphertext_entry =13433205;
#20;
$display("Result = %d", result); assert(result ==6586356);
row = 122;
ciphertext_entry =8678602;
#20;
$display("Result = %d", result); assert(result ==143586);
row = 123;
ciphertext_entry =15433985;
#20;
$display("Result = %d", result); assert(result ==12238596);
row = 124;
ciphertext_entry =5716110;
#20;
$display("Result = %d", result); assert(result ==1341970);
row = 125;
ciphertext_entry =157732;
#20;
$display("Result = %d", result); assert(result ==10222014);
row = 126;
ciphertext_entry =8883810;
#20;
$display("Result = %d", result); assert(result ==9439052);
row = 127;
ciphertext_entry =14103754;
#20;
$display("Result = %d", result); assert(result ==8071470);
row = 128;
ciphertext_entry =5606096;
#20;
$display("Result = %d", result); assert(result ==6722782);
ciphertext_select = 0;
row = 129;
#20;
$display("Result = %d", result); assert(result ==6224554);
row = 130;
#20;
$display("Result = %d", result); assert(result ==16586740);
row = 131;
#20;
$display("Result = %d", result); assert(result ==15423662);
row = 132;
#20;
$display("Result = %d", result); assert(result ==1719904);
row = 133;
#20;
$display("Result = %d", result); assert(result ==8190542);
row = 134;
#20;
$display("Result = %d", result); assert(result ==11338602);
row = 135;
#20;
$display("Result = %d", result); assert(result ==10392892);
row = 136;
#20;
$display("Result = %d", result); assert(result ==9006956);
row = 137;
#20;
$display("Result = %d", result); assert(result ==3292368);
row = 138;
#20;
$display("Result = %d", result); assert(result ==8611648);
row = 139;
#20;
$display("Result = %d", result); assert(result ==7124274);
row = 140;
#20;
$display("Result = %d", result); assert(result ==10436460);
row = 141;
#20;
$display("Result = %d", result); assert(result ==9859874);
row = 142;
#20;
$display("Result = %d", result); assert(result ==10294041);
row = 143;
#20;
$display("Result = %d", result); assert(result ==13022056);
row = 144;
#20;
$display("Result = %d", result); assert(result ==8678417);
row = 145;
#20;
$display("Result = %d", result); assert(result ==7434450);
row = 146;
#20;
$display("Result = %d", result); assert(result ==2154989);
row = 147;
#20;
$display("Result = %d", result); assert(result ==6778639);
row = 148;
#20;
$display("Result = %d", result); assert(result ==12350806);
row = 149;
#20;
$display("Result = %d", result); assert(result ==5061493);
row = 150;
#20;
$display("Result = %d", result); assert(result ==7168203);
row = 151;
#20;
$display("Result = %d", result); assert(result ==7025914);
row = 152;
#20;
$display("Result = %d", result); assert(result ==4449689);
row = 153;
#20;
$display("Result = %d", result); assert(result ==2872604);
row = 154;
#20;
$display("Result = %d", result); assert(result ==12899660);
row = 155;
#20;
$display("Result = %d", result); assert(result ==5692860);
row = 156;
#20;
$display("Result = %d", result); assert(result ==9836967);
row = 157;
#20;
$display("Result = %d", result); assert(result ==15021948);
row = 158;
#20;
$display("Result = %d", result); assert(result ==13821166);
row = 159;
#20;
$display("Result = %d", result); assert(result ==3996274);
row = 160;
#20;
$display("Result = %d", result); assert(result ==14920606);
row = 161;
#20;
$display("Result = %d", result); assert(result ==15540543);
row = 162;
#20;
$display("Result = %d", result); assert(result ==15238076);
row = 163;
#20;
$display("Result = %d", result); assert(result ==11504168);
row = 164;
#20;
$display("Result = %d", result); assert(result ==11967712);
row = 165;
#20;
$display("Result = %d", result); assert(result ==12635672);
row = 166;
#20;
$display("Result = %d", result); assert(result ==14449094);
row = 167;
#20;
$display("Result = %d", result); assert(result ==12243276);
row = 168;
#20;
$display("Result = %d", result); assert(result ==5549106);
row = 169;
#20;
$display("Result = %d", result); assert(result ==3484686);
row = 170;
#20;
$display("Result = %d", result); assert(result ==10697566);
row = 171;
#20;
$display("Result = %d", result); assert(result ==8098055);
row = 172;
#20;
$display("Result = %d", result); assert(result ==9449117);
row = 173;
#20;
$display("Result = %d", result); assert(result ==13053520);
row = 174;
#20;
$display("Result = %d", result); assert(result ==13237191);
row = 175;
#20;
$display("Result = %d", result); assert(result ==9286427);
row = 176;
#20;
$display("Result = %d", result); assert(result ==1223656);
row = 177;
#20;
$display("Result = %d", result); assert(result ==7669603);
row = 178;
#20;
$display("Result = %d", result); assert(result ==6914439);
row = 179;
#20;
$display("Result = %d", result); assert(result ==13608078);
row = 180;
#20;
$display("Result = %d", result); assert(result ==11384996);
row = 181;
#20;
$display("Result = %d", result); assert(result ==14712330);
row = 182;
#20;
$display("Result = %d", result); assert(result ==11011705);
row = 183;
#20;
$display("Result = %d", result); assert(result ==5525258);
row = 184;
#20;
$display("Result = %d", result); assert(result ==3293843);
row = 185;
#20;
$display("Result = %d", result); assert(result ==13787439);
row = 186;
#20;
$display("Result = %d", result); assert(result ==5601184);
row = 187;
#20;
$display("Result = %d", result); assert(result ==7775125);
row = 188;
#20;
$display("Result = %d", result); assert(result ==3462549);
row = 189;
#20;
$display("Result = %d", result); assert(result ==13574767);
row = 190;
#20;
$display("Result = %d", result); assert(result ==1772692);
row = 191;
#20;
$display("Result = %d", result); assert(result ==10503379);
row = 192;
#20;
$display("Result = %d", result); assert(result ==12433105);
row = 193;
#20;
$display("Result = %d", result); assert(result ==3402238);
row = 194;
#20;
$display("Result = %d", result); assert(result ==631394);
row = 195;
#20;
$display("Result = %d", result); assert(result ==14591921);
row = 196;
#20;
$display("Result = %d", result); assert(result ==16445580);
row = 197;
#20;
$display("Result = %d", result); assert(result ==13222457);
row = 198;
#20;
$display("Result = %d", result); assert(result ==12060383);
row = 199;
#20;
$display("Result = %d", result); assert(result ==7062047);
row = 200;
#20;
$display("Result = %d", result); assert(result ==5238742);
row = 201;
#20;
$display("Result = %d", result); assert(result ==9191279);
row = 202;
#20;
$display("Result = %d", result); assert(result ==10731057);
row = 203;
#20;
$display("Result = %d", result); assert(result ==8715503);
row = 204;
#20;
$display("Result = %d", result); assert(result ==15233369);
row = 205;
#20;
$display("Result = %d", result); assert(result ==12087298);
row = 206;
#20;
$display("Result = %d", result); assert(result ==9426270);
row = 207;
#20;
$display("Result = %d", result); assert(result ==15789539);
row = 208;
#20;
$display("Result = %d", result); assert(result ==11671277);
row = 209;
#20;
$display("Result = %d", result); assert(result ==9793926);
row = 210;
#20;
$display("Result = %d", result); assert(result ==12157215);
row = 211;
#20;
$display("Result = %d", result); assert(result ==9845430);
row = 212;
#20;
$display("Result = %d", result); assert(result ==11770655);
row = 213;
#20;
$display("Result = %d", result); assert(result ==855935);
row = 214;
#20;
$display("Result = %d", result); assert(result ==5127519);
row = 215;
#20;
$display("Result = %d", result); assert(result ==1176011);
row = 216;
#20;
$display("Result = %d", result); assert(result ==5853149);
row = 217;
#20;
$display("Result = %d", result); assert(result ==16264309);
row = 218;
#20;
$display("Result = %d", result); assert(result ==5249736);
row = 219;
#20;
$display("Result = %d", result); assert(result ==15243976);
row = 220;
#20;
$display("Result = %d", result); assert(result ==8491791);
row = 221;
#20;
$display("Result = %d", result); assert(result ==11398887);
row = 222;
#20;
$display("Result = %d", result); assert(result ==226590);
row = 223;
#20;
$display("Result = %d", result); assert(result ==607289);
row = 224;
#20;
$display("Result = %d", result); assert(result ==16049783);
row = 225;
#20;
$display("Result = %d", result); assert(result ==16679479);
row = 226;
#20;
$display("Result = %d", result); assert(result ==6654225);
row = 227;
#20;
$display("Result = %d", result); assert(result ==8337118);
row = 228;
#20;
$display("Result = %d", result); assert(result ==11107191);
row = 229;
#20;
$display("Result = %d", result); assert(result ==762143);
row = 230;
#20;
$display("Result = %d", result); assert(result ==15915565);
row = 231;
#20;
$display("Result = %d", result); assert(result ==12323395);
row = 232;
#20;
$display("Result = %d", result); assert(result ==5110909);
row = 233;
#20;
$display("Result = %d", result); assert(result ==16683947);
row = 234;
#20;
$display("Result = %d", result); assert(result ==13559239);
row = 235;
#20;
$display("Result = %d", result); assert(result ==14246191);
row = 236;
#20;
$display("Result = %d", result); assert(result ==6803032);
row = 237;
#20;
$display("Result = %d", result); assert(result ==6111741);
row = 238;
#20;
$display("Result = %d", result); assert(result ==3747897);
row = 239;
#20;
$display("Result = %d", result); assert(result ==10948823);
row = 240;
#20;
$display("Result = %d", result); assert(result ==11668768);
row = 241;
#20;
$display("Result = %d", result); assert(result ==8036192);
row = 242;
#20;
$display("Result = %d", result); assert(result ==12410762);
row = 243;
#20;
$display("Result = %d", result); assert(result ==14972027);
row = 244;
#20;
$display("Result = %d", result); assert(result ==10040478);
row = 245;
#20;
$display("Result = %d", result); assert(result ==2037961);
row = 246;
#20;
$display("Result = %d", result); assert(result ==15114826);
row = 247;
#20;
$display("Result = %d", result); assert(result ==4547071);
row = 248;
#20;
$display("Result = %d", result); assert(result ==11899234);
row = 249;
#20;
$display("Result = %d", result); assert(result ==5820112);
row = 250;
#20;
$display("Result = %d", result); assert(result ==12447446);
row = 251;
#20;
$display("Result = %d", result); assert(result ==7836352);
row = 252;
#20;
$display("Result = %d", result); assert(result ==3809968);
row = 253;
#20;
$display("Result = %d", result); assert(result ==9612844);
row = 254;
#20;
$display("Result = %d", result); assert(result ==10691388);
row = 255;
#20;
$display("Result = %d", result); assert(result ==2021116);
row = 256;
#20;
$display("Result = %d", result); assert(result ==11394784);
en=0;
rst_n=0;
#100;
rst_n=1;
#100;
en=1;
#20;
ciphertext_select = 0;
row = 0;
ciphertext_entry =4810478;
#20;
row = 1;
ciphertext_entry =6346132;
#20;
row = 2;
ciphertext_entry =7107557;
#20;
row = 3;
ciphertext_entry =7645925;
#20;
row = 4;
ciphertext_entry =14800962;
#20;
row = 5;
ciphertext_entry =12339648;
#20;
row = 6;
ciphertext_entry =216637;
#20;
row = 7;
ciphertext_entry =9738200;
#20;
row = 8;
ciphertext_entry =14795173;
#20;
row = 9;
ciphertext_entry =1195151;
#20;
row = 10;
ciphertext_entry =16059388;
#20;
row = 11;
ciphertext_entry =10410615;
#20;
row = 12;
ciphertext_entry =255370;
#20;
row = 13;
ciphertext_entry =2575820;
#20;
row = 14;
ciphertext_entry =16105744;
#20;
row = 15;
ciphertext_entry =15146958;
#20;
row = 16;
ciphertext_entry =10989605;
#20;
row = 17;
ciphertext_entry =6577339;
#20;
row = 18;
ciphertext_entry =8673119;
#20;
row = 19;
ciphertext_entry =10159296;
#20;
row = 20;
ciphertext_entry =12472387;
#20;
row = 21;
ciphertext_entry =16215134;
#20;
row = 22;
ciphertext_entry =212303;
#20;
row = 23;
ciphertext_entry =4878213;
#20;
row = 24;
ciphertext_entry =3160891;
#20;
row = 25;
ciphertext_entry =13441340;
#20;
row = 26;
ciphertext_entry =3824891;
#20;
row = 27;
ciphertext_entry =781959;
#20;
row = 28;
ciphertext_entry =15468565;
#20;
row = 29;
ciphertext_entry =3866432;
#20;
row = 30;
ciphertext_entry =13088017;
#20;
row = 31;
ciphertext_entry =14967363;
#20;
row = 32;
ciphertext_entry =15074930;
#20;
row = 33;
ciphertext_entry =6320442;
#20;
row = 34;
ciphertext_entry =11411877;
#20;
row = 35;
ciphertext_entry =1052583;
#20;
row = 36;
ciphertext_entry =4435825;
#20;
row = 37;
ciphertext_entry =12090247;
#20;
row = 38;
ciphertext_entry =128771;
#20;
row = 39;
ciphertext_entry =15838904;
#20;
row = 40;
ciphertext_entry =10230516;
#20;
row = 41;
ciphertext_entry =5491423;
#20;
row = 42;
ciphertext_entry =7962682;
#20;
row = 43;
ciphertext_entry =9362385;
#20;
row = 44;
ciphertext_entry =8294902;
#20;
row = 45;
ciphertext_entry =4250053;
#20;
row = 46;
ciphertext_entry =13604826;
#20;
row = 47;
ciphertext_entry =9178511;
#20;
row = 48;
ciphertext_entry =6896318;
#20;
row = 49;
ciphertext_entry =6974982;
#20;
row = 50;
ciphertext_entry =1037236;
#20;
row = 51;
ciphertext_entry =431328;
#20;
row = 52;
ciphertext_entry =6909264;
#20;
row = 53;
ciphertext_entry =1877762;
#20;
row = 54;
ciphertext_entry =6259858;
#20;
row = 55;
ciphertext_entry =7436145;
#20;
row = 56;
ciphertext_entry =866009;
#20;
row = 57;
ciphertext_entry =13553724;
#20;
row = 58;
ciphertext_entry =11514901;
#20;
row = 59;
ciphertext_entry =11542027;
#20;
row = 60;
ciphertext_entry =6061506;
#20;
row = 61;
ciphertext_entry =14592150;
#20;
row = 62;
ciphertext_entry =11725663;
#20;
row = 63;
ciphertext_entry =11511778;
#20;
row = 64;
ciphertext_entry =3815008;
#20;
row = 65;
ciphertext_entry =9699081;
#20;
row = 66;
ciphertext_entry =5014095;
#20;
row = 67;
ciphertext_entry =5604246;
#20;
row = 68;
ciphertext_entry =5057791;
#20;
row = 69;
ciphertext_entry =8125737;
#20;
row = 70;
ciphertext_entry =6778074;
#20;
row = 71;
ciphertext_entry =1567253;
#20;
row = 72;
ciphertext_entry =3046989;
#20;
row = 73;
ciphertext_entry =12276548;
#20;
row = 74;
ciphertext_entry =4676664;
#20;
row = 75;
ciphertext_entry =14932871;
#20;
row = 76;
ciphertext_entry =3144818;
#20;
row = 77;
ciphertext_entry =8448975;
#20;
row = 78;
ciphertext_entry =15914698;
#20;
row = 79;
ciphertext_entry =6535121;
#20;
row = 80;
ciphertext_entry =5259203;
#20;
row = 81;
ciphertext_entry =2813274;
#20;
row = 82;
ciphertext_entry =13871045;
#20;
row = 83;
ciphertext_entry =12060141;
#20;
row = 84;
ciphertext_entry =803429;
#20;
row = 85;
ciphertext_entry =7038178;
#20;
row = 86;
ciphertext_entry =11330012;
#20;
row = 87;
ciphertext_entry =4081365;
#20;
row = 88;
ciphertext_entry =661168;
#20;
row = 89;
ciphertext_entry =358866;
#20;
row = 90;
ciphertext_entry =3395483;
#20;
row = 91;
ciphertext_entry =5080712;
#20;
row = 92;
ciphertext_entry =14883804;
#20;
row = 93;
ciphertext_entry =1326218;
#20;
row = 94;
ciphertext_entry =2155744;
#20;
row = 95;
ciphertext_entry =14538235;
#20;
row = 96;
ciphertext_entry =8428683;
#20;
row = 97;
ciphertext_entry =11072099;
#20;
row = 98;
ciphertext_entry =12848853;
#20;
row = 99;
ciphertext_entry =4572389;
#20;
row = 100;
ciphertext_entry =3975828;
#20;
row = 101;
ciphertext_entry =13975293;
#20;
row = 102;
ciphertext_entry =15979760;
#20;
row = 103;
ciphertext_entry =3016031;
#20;
row = 104;
ciphertext_entry =11912223;
#20;
row = 105;
ciphertext_entry =12580149;
#20;
row = 106;
ciphertext_entry =14801902;
#20;
row = 107;
ciphertext_entry =1914548;
#20;
row = 108;
ciphertext_entry =13056952;
#20;
row = 109;
ciphertext_entry =7000225;
#20;
row = 110;
ciphertext_entry =12271218;
#20;
row = 111;
ciphertext_entry =3694931;
#20;
row = 112;
ciphertext_entry =11616085;
#20;
row = 113;
ciphertext_entry =6617547;
#20;
row = 114;
ciphertext_entry =8162162;
#20;
row = 115;
ciphertext_entry =1189603;
#20;
row = 116;
ciphertext_entry =11428240;
#20;
row = 117;
ciphertext_entry =6851109;
#20;
row = 118;
ciphertext_entry =12537811;
#20;
row = 119;
ciphertext_entry =7801557;
#20;
row = 120;
ciphertext_entry =11257284;
#20;
row = 121;
ciphertext_entry =6376319;
#20;
row = 122;
ciphertext_entry =6531035;
#20;
row = 123;
ciphertext_entry =4428540;
#20;
row = 124;
ciphertext_entry =15428460;
#20;
row = 125;
ciphertext_entry =14618815;
#20;
row = 126;
ciphertext_entry =8871752;
#20;
row = 127;
ciphertext_entry =10567613;
#20;
row = 128;
ciphertext_entry =732869;
#20;
ciphertext_select = 1;
row = 0;
ciphertext_entry =4810478;
#20;
$display("Result = %d", result); assert(result ==4686644);
row = 1;
ciphertext_entry =6346132;
#20;
$display("Result = %d", result); assert(result ==4223926);
row = 2;
ciphertext_entry =7107557;
#20;
$display("Result = %d", result); assert(result ==2879416);
row = 3;
ciphertext_entry =7645925;
#20;
$display("Result = %d", result); assert(result ==12186373);
row = 4;
ciphertext_entry =14800962;
#20;
$display("Result = %d", result); assert(result ==15464100);
row = 5;
ciphertext_entry =12339648;
#20;
$display("Result = %d", result); assert(result ==4473240);
row = 6;
ciphertext_entry =216637;
#20;
$display("Result = %d", result); assert(result ==8929476);
row = 7;
ciphertext_entry =9738200;
#20;
$display("Result = %d", result); assert(result ==16138128);
row = 8;
ciphertext_entry =14795173;
#20;
$display("Result = %d", result); assert(result ==4271824);
row = 9;
ciphertext_entry =1195151;
#20;
$display("Result = %d", result); assert(result ==12642791);
row = 10;
ciphertext_entry =16059388;
#20;
$display("Result = %d", result); assert(result ==2352857);
row = 11;
ciphertext_entry =10410615;
#20;
$display("Result = %d", result); assert(result ==3770271);
row = 12;
ciphertext_entry =255370;
#20;
$display("Result = %d", result); assert(result ==6901920);
row = 13;
ciphertext_entry =2575820;
#20;
$display("Result = %d", result); assert(result ==6261999);
row = 14;
ciphertext_entry =16105744;
#20;
$display("Result = %d", result); assert(result ==12232507);
row = 15;
ciphertext_entry =15146958;
#20;
$display("Result = %d", result); assert(result ==8087744);
row = 16;
ciphertext_entry =10989605;
#20;
$display("Result = %d", result); assert(result ==15697108);
row = 17;
ciphertext_entry =6577339;
#20;
$display("Result = %d", result); assert(result ==4808227);
row = 18;
ciphertext_entry =8673119;
#20;
$display("Result = %d", result); assert(result ==11063683);
row = 19;
ciphertext_entry =10159296;
#20;
$display("Result = %d", result); assert(result ==1941768);
row = 20;
ciphertext_entry =12472387;
#20;
$display("Result = %d", result); assert(result ==13472556);
row = 21;
ciphertext_entry =16215134;
#20;
$display("Result = %d", result); assert(result ==9804670);
row = 22;
ciphertext_entry =212303;
#20;
$display("Result = %d", result); assert(result ==11005238);
row = 23;
ciphertext_entry =4878213;
#20;
$display("Result = %d", result); assert(result ==4069885);
row = 24;
ciphertext_entry =3160891;
#20;
$display("Result = %d", result); assert(result ==10734064);
row = 25;
ciphertext_entry =13441340;
#20;
$display("Result = %d", result); assert(result ==470893);
row = 26;
ciphertext_entry =3824891;
#20;
$display("Result = %d", result); assert(result ==2359371);
row = 27;
ciphertext_entry =781959;
#20;
$display("Result = %d", result); assert(result ==13949989);
row = 28;
ciphertext_entry =15468565;
#20;
$display("Result = %d", result); assert(result ==13813910);
row = 29;
ciphertext_entry =3866432;
#20;
$display("Result = %d", result); assert(result ==1057312);
row = 30;
ciphertext_entry =13088017;
#20;
$display("Result = %d", result); assert(result ==10061261);
row = 31;
ciphertext_entry =14967363;
#20;
$display("Result = %d", result); assert(result ==9775208);
row = 32;
ciphertext_entry =15074930;
#20;
$display("Result = %d", result); assert(result ==14375151);
row = 33;
ciphertext_entry =6320442;
#20;
$display("Result = %d", result); assert(result ==694220);
row = 34;
ciphertext_entry =11411877;
#20;
$display("Result = %d", result); assert(result ==7446218);
row = 35;
ciphertext_entry =1052583;
#20;
$display("Result = %d", result); assert(result ==9401463);
row = 36;
ciphertext_entry =4435825;
#20;
$display("Result = %d", result); assert(result ==4782692);
row = 37;
ciphertext_entry =12090247;
#20;
$display("Result = %d", result); assert(result ==15998979);
row = 38;
ciphertext_entry =128771;
#20;
$display("Result = %d", result); assert(result ==10788042);
row = 39;
ciphertext_entry =15838904;
#20;
$display("Result = %d", result); assert(result ==1443585);
row = 40;
ciphertext_entry =10230516;
#20;
$display("Result = %d", result); assert(result ==13373910);
row = 41;
ciphertext_entry =5491423;
#20;
$display("Result = %d", result); assert(result ==13899071);
row = 42;
ciphertext_entry =7962682;
#20;
$display("Result = %d", result); assert(result ==14594810);
row = 43;
ciphertext_entry =9362385;
#20;
$display("Result = %d", result); assert(result ==9771842);
row = 44;
ciphertext_entry =8294902;
#20;
$display("Result = %d", result); assert(result ==8874829);
row = 45;
ciphertext_entry =4250053;
#20;
$display("Result = %d", result); assert(result ==7036621);
row = 46;
ciphertext_entry =13604826;
#20;
$display("Result = %d", result); assert(result ==7381916);
row = 47;
ciphertext_entry =9178511;
#20;
$display("Result = %d", result); assert(result ==8822470);
row = 48;
ciphertext_entry =6896318;
#20;
$display("Result = %d", result); assert(result ==16352068);
row = 49;
ciphertext_entry =6974982;
#20;
$display("Result = %d", result); assert(result ==11946334);
row = 50;
ciphertext_entry =1037236;
#20;
$display("Result = %d", result); assert(result ==8046107);
row = 51;
ciphertext_entry =431328;
#20;
$display("Result = %d", result); assert(result ==10186456);
row = 52;
ciphertext_entry =6909264;
#20;
$display("Result = %d", result); assert(result ==742352);
row = 53;
ciphertext_entry =1877762;
#20;
$display("Result = %d", result); assert(result ==3111139);
row = 54;
ciphertext_entry =6259858;
#20;
$display("Result = %d", result); assert(result ==5577107);
row = 55;
ciphertext_entry =7436145;
#20;
$display("Result = %d", result); assert(result ==11522451);
row = 56;
ciphertext_entry =866009;
#20;
$display("Result = %d", result); assert(result ==11639387);
row = 57;
ciphertext_entry =13553724;
#20;
$display("Result = %d", result); assert(result ==8532414);
row = 58;
ciphertext_entry =11514901;
#20;
$display("Result = %d", result); assert(result ==2370578);
row = 59;
ciphertext_entry =11542027;
#20;
$display("Result = %d", result); assert(result ==7233256);
row = 60;
ciphertext_entry =6061506;
#20;
$display("Result = %d", result); assert(result ==7954875);
row = 61;
ciphertext_entry =14592150;
#20;
$display("Result = %d", result); assert(result ==3452439);
row = 62;
ciphertext_entry =11725663;
#20;
$display("Result = %d", result); assert(result ==6329023);
row = 63;
ciphertext_entry =11511778;
#20;
$display("Result = %d", result); assert(result ==3898685);
row = 64;
ciphertext_entry =3815008;
#20;
$display("Result = %d", result); assert(result ==13246130);
row = 65;
ciphertext_entry =9699081;
#20;
$display("Result = %d", result); assert(result ==7258255);
row = 66;
ciphertext_entry =5014095;
#20;
$display("Result = %d", result); assert(result ==15680840);
row = 67;
ciphertext_entry =5604246;
#20;
$display("Result = %d", result); assert(result ==3482221);
row = 68;
ciphertext_entry =5057791;
#20;
$display("Result = %d", result); assert(result ==7576629);
row = 69;
ciphertext_entry =8125737;
#20;
$display("Result = %d", result); assert(result ==6738756);
row = 70;
ciphertext_entry =6778074;
#20;
$display("Result = %d", result); assert(result ==547121);
row = 71;
ciphertext_entry =1567253;
#20;
$display("Result = %d", result); assert(result ==16554624);
row = 72;
ciphertext_entry =3046989;
#20;
$display("Result = %d", result); assert(result ==12863415);
row = 73;
ciphertext_entry =12276548;
#20;
$display("Result = %d", result); assert(result ==11117132);
row = 74;
ciphertext_entry =4676664;
#20;
$display("Result = %d", result); assert(result ==6633172);
row = 75;
ciphertext_entry =14932871;
#20;
$display("Result = %d", result); assert(result ==6158287);
row = 76;
ciphertext_entry =3144818;
#20;
$display("Result = %d", result); assert(result ==5035534);
row = 77;
ciphertext_entry =8448975;
#20;
$display("Result = %d", result); assert(result ==2307547);
row = 78;
ciphertext_entry =15914698;
#20;
$display("Result = %d", result); assert(result ==2717396);
row = 79;
ciphertext_entry =6535121;
#20;
$display("Result = %d", result); assert(result ==4088169);
row = 80;
ciphertext_entry =5259203;
#20;
$display("Result = %d", result); assert(result ==17586);
row = 81;
ciphertext_entry =2813274;
#20;
$display("Result = %d", result); assert(result ==3105402);
row = 82;
ciphertext_entry =13871045;
#20;
$display("Result = %d", result); assert(result ==10686288);
row = 83;
ciphertext_entry =12060141;
#20;
$display("Result = %d", result); assert(result ==16483821);
row = 84;
ciphertext_entry =803429;
#20;
$display("Result = %d", result); assert(result ==10390560);
row = 85;
ciphertext_entry =7038178;
#20;
$display("Result = %d", result); assert(result ==13665512);
row = 86;
ciphertext_entry =11330012;
#20;
$display("Result = %d", result); assert(result ==1039509);
row = 87;
ciphertext_entry =4081365;
#20;
$display("Result = %d", result); assert(result ==9488635);
row = 88;
ciphertext_entry =661168;
#20;
$display("Result = %d", result); assert(result ==7256628);
row = 89;
ciphertext_entry =358866;
#20;
$display("Result = %d", result); assert(result ==11874904);
row = 90;
ciphertext_entry =3395483;
#20;
$display("Result = %d", result); assert(result ==3940829);
row = 91;
ciphertext_entry =5080712;
#20;
$display("Result = %d", result); assert(result ==1669057);
row = 92;
ciphertext_entry =14883804;
#20;
$display("Result = %d", result); assert(result ==1701644);
row = 93;
ciphertext_entry =1326218;
#20;
$display("Result = %d", result); assert(result ==6990475);
row = 94;
ciphertext_entry =2155744;
#20;
$display("Result = %d", result); assert(result ==11873009);
row = 95;
ciphertext_entry =14538235;
#20;
$display("Result = %d", result); assert(result ==16221944);
row = 96;
ciphertext_entry =8428683;
#20;
$display("Result = %d", result); assert(result ==3782199);
row = 97;
ciphertext_entry =11072099;
#20;
$display("Result = %d", result); assert(result ==7164250);
row = 98;
ciphertext_entry =12848853;
#20;
$display("Result = %d", result); assert(result ==4272719);
row = 99;
ciphertext_entry =4572389;
#20;
$display("Result = %d", result); assert(result ==10129692);
row = 100;
ciphertext_entry =3975828;
#20;
$display("Result = %d", result); assert(result ==1333700);
row = 101;
ciphertext_entry =13975293;
#20;
$display("Result = %d", result); assert(result ==12768188);
row = 102;
ciphertext_entry =15979760;
#20;
$display("Result = %d", result); assert(result ==3641309);
row = 103;
ciphertext_entry =3016031;
#20;
$display("Result = %d", result); assert(result ==11671050);
row = 104;
ciphertext_entry =11912223;
#20;
$display("Result = %d", result); assert(result ==9585189);
row = 105;
ciphertext_entry =12580149;
#20;
$display("Result = %d", result); assert(result ==7953542);
row = 106;
ciphertext_entry =14801902;
#20;
$display("Result = %d", result); assert(result ==6489742);
row = 107;
ciphertext_entry =1914548;
#20;
$display("Result = %d", result); assert(result ==9459855);
row = 108;
ciphertext_entry =13056952;
#20;
$display("Result = %d", result); assert(result ==7473637);
row = 109;
ciphertext_entry =7000225;
#20;
$display("Result = %d", result); assert(result ==2591381);
row = 110;
ciphertext_entry =12271218;
#20;
$display("Result = %d", result); assert(result ==8763380);
row = 111;
ciphertext_entry =3694931;
#20;
$display("Result = %d", result); assert(result ==9265672);
row = 112;
ciphertext_entry =11616085;
#20;
$display("Result = %d", result); assert(result ==7826361);
row = 113;
ciphertext_entry =6617547;
#20;
$display("Result = %d", result); assert(result ==7356562);
row = 114;
ciphertext_entry =8162162;
#20;
$display("Result = %d", result); assert(result ==2625069);
row = 115;
ciphertext_entry =1189603;
#20;
$display("Result = %d", result); assert(result ==10694789);
row = 116;
ciphertext_entry =11428240;
#20;
$display("Result = %d", result); assert(result ==12353858);
row = 117;
ciphertext_entry =6851109;
#20;
$display("Result = %d", result); assert(result ==10427491);
row = 118;
ciphertext_entry =12537811;
#20;
$display("Result = %d", result); assert(result ==13411463);
row = 119;
ciphertext_entry =7801557;
#20;
$display("Result = %d", result); assert(result ==7240169);
row = 120;
ciphertext_entry =11257284;
#20;
$display("Result = %d", result); assert(result ==11409835);
row = 121;
ciphertext_entry =6376319;
#20;
$display("Result = %d", result); assert(result ==6608914);
row = 122;
ciphertext_entry =6531035;
#20;
$display("Result = %d", result); assert(result ==1846632);
row = 123;
ciphertext_entry =4428540;
#20;
$display("Result = %d", result); assert(result ==15094254);
row = 124;
ciphertext_entry =15428460;
#20;
$display("Result = %d", result); assert(result ==4466233);
row = 125;
ciphertext_entry =14618815;
#20;
$display("Result = %d", result); assert(result ==997180);
row = 126;
ciphertext_entry =8871752;
#20;
$display("Result = %d", result); assert(result ==5295508);
row = 127;
ciphertext_entry =10567613;
#20;
$display("Result = %d", result); assert(result ==8881028);
row = 128;
ciphertext_entry =732869;
#20;
$display("Result = %d", result); assert(result ==818789);
ciphertext_select = 0;
row = 129;
#20;
$display("Result = %d", result); assert(result ==2340988);
row = 130;
#20;
$display("Result = %d", result); assert(result ==5774661);
row = 131;
#20;
$display("Result = %d", result); assert(result ==7062074);
row = 132;
#20;
$display("Result = %d", result); assert(result ==3250072);
row = 133;
#20;
$display("Result = %d", result); assert(result ==16190447);
row = 134;
#20;
$display("Result = %d", result); assert(result ==5231674);
row = 135;
#20;
$display("Result = %d", result); assert(result ==3987194);
row = 136;
#20;
$display("Result = %d", result); assert(result ==9551443);
row = 137;
#20;
$display("Result = %d", result); assert(result ==11860317);
row = 138;
#20;
$display("Result = %d", result); assert(result ==13941119);
row = 139;
#20;
$display("Result = %d", result); assert(result ==3278517);
row = 140;
#20;
$display("Result = %d", result); assert(result ==6831238);
row = 141;
#20;
$display("Result = %d", result); assert(result ==9771659);
row = 142;
#20;
$display("Result = %d", result); assert(result ==11150646);
row = 143;
#20;
$display("Result = %d", result); assert(result ==12886725);
row = 144;
#20;
$display("Result = %d", result); assert(result ==9248600);
row = 145;
#20;
$display("Result = %d", result); assert(result ==13120807);
row = 146;
#20;
$display("Result = %d", result); assert(result ==12402722);
row = 147;
#20;
$display("Result = %d", result); assert(result ==1508277);
row = 148;
#20;
$display("Result = %d", result); assert(result ==11983302);
row = 149;
#20;
$display("Result = %d", result); assert(result ==15100211);
row = 150;
#20;
$display("Result = %d", result); assert(result ==7775380);
row = 151;
#20;
$display("Result = %d", result); assert(result ==16075538);
row = 152;
#20;
$display("Result = %d", result); assert(result ==5279255);
row = 153;
#20;
$display("Result = %d", result); assert(result ==1266760);
row = 154;
#20;
$display("Result = %d", result); assert(result ==9092974);
row = 155;
#20;
$display("Result = %d", result); assert(result ==11283530);
row = 156;
#20;
$display("Result = %d", result); assert(result ==953964);
row = 157;
#20;
$display("Result = %d", result); assert(result ==12722373);
row = 158;
#20;
$display("Result = %d", result); assert(result ==11401194);
row = 159;
#20;
$display("Result = %d", result); assert(result ==13461177);
row = 160;
#20;
$display("Result = %d", result); assert(result ==14838632);
row = 161;
#20;
$display("Result = %d", result); assert(result ==6757523);
row = 162;
#20;
$display("Result = %d", result); assert(result ==2739533);
row = 163;
#20;
$display("Result = %d", result); assert(result ==12775450);
row = 164;
#20;
$display("Result = %d", result); assert(result ==12529566);
row = 165;
#20;
$display("Result = %d", result); assert(result ==6132778);
row = 166;
#20;
$display("Result = %d", result); assert(result ==13103783);
row = 167;
#20;
$display("Result = %d", result); assert(result ==363778);
row = 168;
#20;
$display("Result = %d", result); assert(result ==5395925);
row = 169;
#20;
$display("Result = %d", result); assert(result ==8914301);
row = 170;
#20;
$display("Result = %d", result); assert(result ==2618854);
row = 171;
#20;
$display("Result = %d", result); assert(result ==11555894);
row = 172;
#20;
$display("Result = %d", result); assert(result ==14676618);
row = 173;
#20;
$display("Result = %d", result); assert(result ==12421643);
row = 174;
#20;
$display("Result = %d", result); assert(result ==6028177);
row = 175;
#20;
$display("Result = %d", result); assert(result ==14374757);
row = 176;
#20;
$display("Result = %d", result); assert(result ==9140261);
row = 177;
#20;
$display("Result = %d", result); assert(result ==961089);
row = 178;
#20;
$display("Result = %d", result); assert(result ==16744616);
row = 179;
#20;
$display("Result = %d", result); assert(result ==1651284);
row = 180;
#20;
$display("Result = %d", result); assert(result ==12093009);
row = 181;
#20;
$display("Result = %d", result); assert(result ==1575866);
row = 182;
#20;
$display("Result = %d", result); assert(result ==7529764);
row = 183;
#20;
$display("Result = %d", result); assert(result ==15559937);
row = 184;
#20;
$display("Result = %d", result); assert(result ==12764426);
row = 185;
#20;
$display("Result = %d", result); assert(result ==4008396);
row = 186;
#20;
$display("Result = %d", result); assert(result ==8301217);
row = 187;
#20;
$display("Result = %d", result); assert(result ==6155194);
row = 188;
#20;
$display("Result = %d", result); assert(result ==2293579);
row = 189;
#20;
$display("Result = %d", result); assert(result ==8594647);
row = 190;
#20;
$display("Result = %d", result); assert(result ==1069501);
row = 191;
#20;
$display("Result = %d", result); assert(result ==4423333);
row = 192;
#20;
$display("Result = %d", result); assert(result ==427844);
row = 193;
#20;
$display("Result = %d", result); assert(result ==8408410);
row = 194;
#20;
$display("Result = %d", result); assert(result ==7929445);
row = 195;
#20;
$display("Result = %d", result); assert(result ==9672650);
row = 196;
#20;
$display("Result = %d", result); assert(result ==10666540);
row = 197;
#20;
$display("Result = %d", result); assert(result ==12375899);
row = 198;
#20;
$display("Result = %d", result); assert(result ==1557569);
row = 199;
#20;
$display("Result = %d", result); assert(result ==1532374);
row = 200;
#20;
$display("Result = %d", result); assert(result ==6644952);
row = 201;
#20;
$display("Result = %d", result); assert(result ==14917177);
row = 202;
#20;
$display("Result = %d", result); assert(result ==7432798);
row = 203;
#20;
$display("Result = %d", result); assert(result ==5147912);
row = 204;
#20;
$display("Result = %d", result); assert(result ==2810912);
row = 205;
#20;
$display("Result = %d", result); assert(result ==3459424);
row = 206;
#20;
$display("Result = %d", result); assert(result ==7653558);
row = 207;
#20;
$display("Result = %d", result); assert(result ==13587517);
row = 208;
#20;
$display("Result = %d", result); assert(result ==4574496);
row = 209;
#20;
$display("Result = %d", result); assert(result ==5916558);
row = 210;
#20;
$display("Result = %d", result); assert(result ==5654811);
row = 211;
#20;
$display("Result = %d", result); assert(result ==13608104);
row = 212;
#20;
$display("Result = %d", result); assert(result ==14834951);
row = 213;
#20;
$display("Result = %d", result); assert(result ==11760918);
row = 214;
#20;
$display("Result = %d", result); assert(result ==14987649);
row = 215;
#20;
$display("Result = %d", result); assert(result ==3204869);
row = 216;
#20;
$display("Result = %d", result); assert(result ==8900493);
row = 217;
#20;
$display("Result = %d", result); assert(result ==7489982);
row = 218;
#20;
$display("Result = %d", result); assert(result ==9383108);
row = 219;
#20;
$display("Result = %d", result); assert(result ==6431542);
row = 220;
#20;
$display("Result = %d", result); assert(result ==16057059);
row = 221;
#20;
$display("Result = %d", result); assert(result ==3380040);
row = 222;
#20;
$display("Result = %d", result); assert(result ==2701568);
row = 223;
#20;
$display("Result = %d", result); assert(result ==13623845);
row = 224;
#20;
$display("Result = %d", result); assert(result ==1264306);
row = 225;
#20;
$display("Result = %d", result); assert(result ==14511644);
row = 226;
#20;
$display("Result = %d", result); assert(result ==5326528);
row = 227;
#20;
$display("Result = %d", result); assert(result ==15503221);
row = 228;
#20;
$display("Result = %d", result); assert(result ==6867095);
row = 229;
#20;
$display("Result = %d", result); assert(result ==3736205);
row = 230;
#20;
$display("Result = %d", result); assert(result ==15647628);
row = 231;
#20;
$display("Result = %d", result); assert(result ==5983688);
row = 232;
#20;
$display("Result = %d", result); assert(result ==1536653);
row = 233;
#20;
$display("Result = %d", result); assert(result ==15329711);
row = 234;
#20;
$display("Result = %d", result); assert(result ==7569858);
row = 235;
#20;
$display("Result = %d", result); assert(result ==8038127);
row = 236;
#20;
$display("Result = %d", result); assert(result ==5935208);
row = 237;
#20;
$display("Result = %d", result); assert(result ==11993264);
row = 238;
#20;
$display("Result = %d", result); assert(result ==4227719);
row = 239;
#20;
$display("Result = %d", result); assert(result ==2220657);
row = 240;
#20;
$display("Result = %d", result); assert(result ==11244386);
row = 241;
#20;
$display("Result = %d", result); assert(result ==5783863);
row = 242;
#20;
$display("Result = %d", result); assert(result ==16184372);
row = 243;
#20;
$display("Result = %d", result); assert(result ==4552881);
row = 244;
#20;
$display("Result = %d", result); assert(result ==4523315);
row = 245;
#20;
$display("Result = %d", result); assert(result ==4534095);
row = 246;
#20;
$display("Result = %d", result); assert(result ==9817477);
row = 247;
#20;
$display("Result = %d", result); assert(result ==3313214);
row = 248;
#20;
$display("Result = %d", result); assert(result ==2051710);
row = 249;
#20;
$display("Result = %d", result); assert(result ==9230932);
row = 250;
#20;
$display("Result = %d", result); assert(result ==2029267);
row = 251;
#20;
$display("Result = %d", result); assert(result ==3898904);
row = 252;
#20;
$display("Result = %d", result); assert(result ==8494398);
row = 253;
#20;
$display("Result = %d", result); assert(result ==5605358);
row = 254;
#20;
$display("Result = %d", result); assert(result ==5414982);
row = 255;
#20;
$display("Result = %d", result); assert(result ==11610476);
row = 256;
#20;
$display("Result = %d", result); assert(result ==8344916);
en=0;
rst_n=0;
#100;
rst_n=1;
#100;
en=1;
#20;
ciphertext_select = 0;
row = 0;
ciphertext_entry =7065155;
#20;
row = 1;
ciphertext_entry =7210534;
#20;
row = 2;
ciphertext_entry =4818605;
#20;
row = 3;
ciphertext_entry =1138268;
#20;
row = 4;
ciphertext_entry =14366918;
#20;
row = 5;
ciphertext_entry =11700516;
#20;
row = 6;
ciphertext_entry =10008479;
#20;
row = 7;
ciphertext_entry =10466143;
#20;
row = 8;
ciphertext_entry =6428024;
#20;
row = 9;
ciphertext_entry =5394108;
#20;
row = 10;
ciphertext_entry =2718485;
#20;
row = 11;
ciphertext_entry =12088624;
#20;
row = 12;
ciphertext_entry =16149648;
#20;
row = 13;
ciphertext_entry =309070;
#20;
row = 14;
ciphertext_entry =6368466;
#20;
row = 15;
ciphertext_entry =16739327;
#20;
row = 16;
ciphertext_entry =2416418;
#20;
row = 17;
ciphertext_entry =12361961;
#20;
row = 18;
ciphertext_entry =8715868;
#20;
row = 19;
ciphertext_entry =10451330;
#20;
row = 20;
ciphertext_entry =12117999;
#20;
row = 21;
ciphertext_entry =5486688;
#20;
row = 22;
ciphertext_entry =8159486;
#20;
row = 23;
ciphertext_entry =15809805;
#20;
row = 24;
ciphertext_entry =13746083;
#20;
row = 25;
ciphertext_entry =1548111;
#20;
row = 26;
ciphertext_entry =11387475;
#20;
row = 27;
ciphertext_entry =4024491;
#20;
row = 28;
ciphertext_entry =13807856;
#20;
row = 29;
ciphertext_entry =12660493;
#20;
row = 30;
ciphertext_entry =14421618;
#20;
row = 31;
ciphertext_entry =5516472;
#20;
row = 32;
ciphertext_entry =10753472;
#20;
row = 33;
ciphertext_entry =14923305;
#20;
row = 34;
ciphertext_entry =11276310;
#20;
row = 35;
ciphertext_entry =4119004;
#20;
row = 36;
ciphertext_entry =2220252;
#20;
row = 37;
ciphertext_entry =15422095;
#20;
row = 38;
ciphertext_entry =13964385;
#20;
row = 39;
ciphertext_entry =7440141;
#20;
row = 40;
ciphertext_entry =8189649;
#20;
row = 41;
ciphertext_entry =3381218;
#20;
row = 42;
ciphertext_entry =3720981;
#20;
row = 43;
ciphertext_entry =318102;
#20;
row = 44;
ciphertext_entry =4412987;
#20;
row = 45;
ciphertext_entry =3746988;
#20;
row = 46;
ciphertext_entry =2967712;
#20;
row = 47;
ciphertext_entry =5765138;
#20;
row = 48;
ciphertext_entry =2997420;
#20;
row = 49;
ciphertext_entry =9642920;
#20;
row = 50;
ciphertext_entry =16723935;
#20;
row = 51;
ciphertext_entry =16183603;
#20;
row = 52;
ciphertext_entry =15017472;
#20;
row = 53;
ciphertext_entry =13782877;
#20;
row = 54;
ciphertext_entry =2886937;
#20;
row = 55;
ciphertext_entry =12764177;
#20;
row = 56;
ciphertext_entry =9979893;
#20;
row = 57;
ciphertext_entry =9714129;
#20;
row = 58;
ciphertext_entry =10696438;
#20;
row = 59;
ciphertext_entry =14360916;
#20;
row = 60;
ciphertext_entry =8337423;
#20;
row = 61;
ciphertext_entry =2247231;
#20;
row = 62;
ciphertext_entry =8277517;
#20;
row = 63;
ciphertext_entry =10964515;
#20;
row = 64;
ciphertext_entry =9290115;
#20;
row = 65;
ciphertext_entry =15266607;
#20;
row = 66;
ciphertext_entry =8902809;
#20;
row = 67;
ciphertext_entry =7897649;
#20;
row = 68;
ciphertext_entry =10773300;
#20;
row = 69;
ciphertext_entry =11945652;
#20;
row = 70;
ciphertext_entry =7475770;
#20;
row = 71;
ciphertext_entry =6464462;
#20;
row = 72;
ciphertext_entry =8445158;
#20;
row = 73;
ciphertext_entry =11422268;
#20;
row = 74;
ciphertext_entry =15171220;
#20;
row = 75;
ciphertext_entry =598323;
#20;
row = 76;
ciphertext_entry =12282367;
#20;
row = 77;
ciphertext_entry =9312931;
#20;
row = 78;
ciphertext_entry =5802789;
#20;
row = 79;
ciphertext_entry =8048348;
#20;
row = 80;
ciphertext_entry =2613732;
#20;
row = 81;
ciphertext_entry =13810549;
#20;
row = 82;
ciphertext_entry =1025754;
#20;
row = 83;
ciphertext_entry =1300761;
#20;
row = 84;
ciphertext_entry =14396277;
#20;
row = 85;
ciphertext_entry =13247639;
#20;
row = 86;
ciphertext_entry =7378534;
#20;
row = 87;
ciphertext_entry =13578534;
#20;
row = 88;
ciphertext_entry =6631803;
#20;
row = 89;
ciphertext_entry =6539247;
#20;
row = 90;
ciphertext_entry =9670700;
#20;
row = 91;
ciphertext_entry =12541800;
#20;
row = 92;
ciphertext_entry =662742;
#20;
row = 93;
ciphertext_entry =14810215;
#20;
row = 94;
ciphertext_entry =14564306;
#20;
row = 95;
ciphertext_entry =15812604;
#20;
row = 96;
ciphertext_entry =878920;
#20;
row = 97;
ciphertext_entry =1179072;
#20;
row = 98;
ciphertext_entry =11098319;
#20;
row = 99;
ciphertext_entry =6504697;
#20;
row = 100;
ciphertext_entry =5157978;
#20;
row = 101;
ciphertext_entry =6349629;
#20;
row = 102;
ciphertext_entry =3513589;
#20;
row = 103;
ciphertext_entry =9104225;
#20;
row = 104;
ciphertext_entry =14514092;
#20;
row = 105;
ciphertext_entry =435730;
#20;
row = 106;
ciphertext_entry =3124935;
#20;
row = 107;
ciphertext_entry =7082632;
#20;
row = 108;
ciphertext_entry =15306750;
#20;
row = 109;
ciphertext_entry =10252241;
#20;
row = 110;
ciphertext_entry =1517219;
#20;
row = 111;
ciphertext_entry =12865329;
#20;
row = 112;
ciphertext_entry =6884282;
#20;
row = 113;
ciphertext_entry =16527876;
#20;
row = 114;
ciphertext_entry =4831239;
#20;
row = 115;
ciphertext_entry =13777612;
#20;
row = 116;
ciphertext_entry =9520487;
#20;
row = 117;
ciphertext_entry =1068946;
#20;
row = 118;
ciphertext_entry =1295344;
#20;
row = 119;
ciphertext_entry =14240044;
#20;
row = 120;
ciphertext_entry =11943159;
#20;
row = 121;
ciphertext_entry =8016467;
#20;
row = 122;
ciphertext_entry =9559681;
#20;
row = 123;
ciphertext_entry =3361994;
#20;
row = 124;
ciphertext_entry =3826283;
#20;
row = 125;
ciphertext_entry =16026884;
#20;
row = 126;
ciphertext_entry =15484096;
#20;
row = 127;
ciphertext_entry =562818;
#20;
row = 128;
ciphertext_entry =13170074;
#20;
ciphertext_select = 1;
row = 0;
ciphertext_entry =7065155;
#20;
$display("Result = %d", result); assert(result ==15137702);
row = 1;
ciphertext_entry =7210534;
#20;
$display("Result = %d", result); assert(result ==15498276);
row = 2;
ciphertext_entry =4818605;
#20;
$display("Result = %d", result); assert(result ==10450869);
row = 3;
ciphertext_entry =1138268;
#20;
$display("Result = %d", result); assert(result ==13970119);
row = 4;
ciphertext_entry =14366918;
#20;
$display("Result = %d", result); assert(result ==3922410);
row = 5;
ciphertext_entry =11700516;
#20;
$display("Result = %d", result); assert(result ==11863757);
row = 6;
ciphertext_entry =10008479;
#20;
$display("Result = %d", result); assert(result ==5367131);
row = 7;
ciphertext_entry =10466143;
#20;
$display("Result = %d", result); assert(result ==16649298);
row = 8;
ciphertext_entry =6428024;
#20;
$display("Result = %d", result); assert(result ==4548081);
row = 9;
ciphertext_entry =5394108;
#20;
$display("Result = %d", result); assert(result ==123244);
row = 10;
ciphertext_entry =2718485;
#20;
$display("Result = %d", result); assert(result ==13691328);
row = 11;
ciphertext_entry =12088624;
#20;
$display("Result = %d", result); assert(result ==1645113);
row = 12;
ciphertext_entry =16149648;
#20;
$display("Result = %d", result); assert(result ==8731085);
row = 13;
ciphertext_entry =309070;
#20;
$display("Result = %d", result); assert(result ==6707454);
row = 14;
ciphertext_entry =6368466;
#20;
$display("Result = %d", result); assert(result ==12180953);
row = 15;
ciphertext_entry =16739327;
#20;
$display("Result = %d", result); assert(result ==692674);
row = 16;
ciphertext_entry =2416418;
#20;
$display("Result = %d", result); assert(result ==10864757);
row = 17;
ciphertext_entry =12361961;
#20;
$display("Result = %d", result); assert(result ==15839739);
row = 18;
ciphertext_entry =8715868;
#20;
$display("Result = %d", result); assert(result ==13025151);
row = 19;
ciphertext_entry =10451330;
#20;
$display("Result = %d", result); assert(result ==11762734);
row = 20;
ciphertext_entry =12117999;
#20;
$display("Result = %d", result); assert(result ==7580319);
row = 21;
ciphertext_entry =5486688;
#20;
$display("Result = %d", result); assert(result ==7323456);
row = 22;
ciphertext_entry =8159486;
#20;
$display("Result = %d", result); assert(result ==13540558);
row = 23;
ciphertext_entry =15809805;
#20;
$display("Result = %d", result); assert(result ==9505588);
row = 24;
ciphertext_entry =13746083;
#20;
$display("Result = %d", result); assert(result ==11512641);
row = 25;
ciphertext_entry =1548111;
#20;
$display("Result = %d", result); assert(result ==16398323);
row = 26;
ciphertext_entry =11387475;
#20;
$display("Result = %d", result); assert(result ==2627506);
row = 27;
ciphertext_entry =4024491;
#20;
$display("Result = %d", result); assert(result ==9709537);
row = 28;
ciphertext_entry =13807856;
#20;
$display("Result = %d", result); assert(result ==16136153);
row = 29;
ciphertext_entry =12660493;
#20;
$display("Result = %d", result); assert(result ==14068490);
row = 30;
ciphertext_entry =14421618;
#20;
$display("Result = %d", result); assert(result ==9439862);
row = 31;
ciphertext_entry =5516472;
#20;
$display("Result = %d", result); assert(result ==7695468);
row = 32;
ciphertext_entry =10753472;
#20;
$display("Result = %d", result); assert(result ==15286714);
row = 33;
ciphertext_entry =14923305;
#20;
$display("Result = %d", result); assert(result ==1068220);
row = 34;
ciphertext_entry =11276310;
#20;
$display("Result = %d", result); assert(result ==7396116);
row = 35;
ciphertext_entry =4119004;
#20;
$display("Result = %d", result); assert(result ==13799982);
row = 36;
ciphertext_entry =2220252;
#20;
$display("Result = %d", result); assert(result ==2040981);
row = 37;
ciphertext_entry =15422095;
#20;
$display("Result = %d", result); assert(result ==13380646);
row = 38;
ciphertext_entry =13964385;
#20;
$display("Result = %d", result); assert(result ==6405457);
row = 39;
ciphertext_entry =7440141;
#20;
$display("Result = %d", result); assert(result ==10886336);
row = 40;
ciphertext_entry =8189649;
#20;
$display("Result = %d", result); assert(result ==8996093);
row = 41;
ciphertext_entry =3381218;
#20;
$display("Result = %d", result); assert(result ==7786443);
row = 42;
ciphertext_entry =3720981;
#20;
$display("Result = %d", result); assert(result ==5189486);
row = 43;
ciphertext_entry =318102;
#20;
$display("Result = %d", result); assert(result ==13405531);
row = 44;
ciphertext_entry =4412987;
#20;
$display("Result = %d", result); assert(result ==13636326);
row = 45;
ciphertext_entry =3746988;
#20;
$display("Result = %d", result); assert(result ==12573671);
row = 46;
ciphertext_entry =2967712;
#20;
$display("Result = %d", result); assert(result ==6180993);
row = 47;
ciphertext_entry =5765138;
#20;
$display("Result = %d", result); assert(result ==13208668);
row = 48;
ciphertext_entry =2997420;
#20;
$display("Result = %d", result); assert(result ==9477456);
row = 49;
ciphertext_entry =9642920;
#20;
$display("Result = %d", result); assert(result ==1187504);
row = 50;
ciphertext_entry =16723935;
#20;
$display("Result = %d", result); assert(result ==7576107);
row = 51;
ciphertext_entry =16183603;
#20;
$display("Result = %d", result); assert(result ==13004128);
row = 52;
ciphertext_entry =15017472;
#20;
$display("Result = %d", result); assert(result ==2770603);
row = 53;
ciphertext_entry =13782877;
#20;
$display("Result = %d", result); assert(result ==6206713);
row = 54;
ciphertext_entry =2886937;
#20;
$display("Result = %d", result); assert(result ==12088793);
row = 55;
ciphertext_entry =12764177;
#20;
$display("Result = %d", result); assert(result ==16649893);
row = 56;
ciphertext_entry =9979893;
#20;
$display("Result = %d", result); assert(result ==12771387);
row = 57;
ciphertext_entry =9714129;
#20;
$display("Result = %d", result); assert(result ==2242244);
row = 58;
ciphertext_entry =10696438;
#20;
$display("Result = %d", result); assert(result ==10825929);
row = 59;
ciphertext_entry =14360916;
#20;
$display("Result = %d", result); assert(result ==10598402);
row = 60;
ciphertext_entry =8337423;
#20;
$display("Result = %d", result); assert(result ==4456459);
row = 61;
ciphertext_entry =2247231;
#20;
$display("Result = %d", result); assert(result ==9779550);
row = 62;
ciphertext_entry =8277517;
#20;
$display("Result = %d", result); assert(result ==5619123);
row = 63;
ciphertext_entry =10964515;
#20;
$display("Result = %d", result); assert(result ==3822221);
row = 64;
ciphertext_entry =9290115;
#20;
$display("Result = %d", result); assert(result ==14325305);
row = 65;
ciphertext_entry =15266607;
#20;
$display("Result = %d", result); assert(result ==5436524);
row = 66;
ciphertext_entry =8902809;
#20;
$display("Result = %d", result); assert(result ==10567649);
row = 67;
ciphertext_entry =7897649;
#20;
$display("Result = %d", result); assert(result ==5774443);
row = 68;
ciphertext_entry =10773300;
#20;
$display("Result = %d", result); assert(result ==16193207);
row = 69;
ciphertext_entry =11945652;
#20;
$display("Result = %d", result); assert(result ==11901481);
row = 70;
ciphertext_entry =7475770;
#20;
$display("Result = %d", result); assert(result ==1514930);
row = 71;
ciphertext_entry =6464462;
#20;
$display("Result = %d", result); assert(result ==7650931);
row = 72;
ciphertext_entry =8445158;
#20;
$display("Result = %d", result); assert(result ==16475093);
row = 73;
ciphertext_entry =11422268;
#20;
$display("Result = %d", result); assert(result ==14755442);
row = 74;
ciphertext_entry =15171220;
#20;
$display("Result = %d", result); assert(result ==335598);
row = 75;
ciphertext_entry =598323;
#20;
$display("Result = %d", result); assert(result ==5086192);
row = 76;
ciphertext_entry =12282367;
#20;
$display("Result = %d", result); assert(result ==16095541);
row = 77;
ciphertext_entry =9312931;
#20;
$display("Result = %d", result); assert(result ==1189144);
row = 78;
ciphertext_entry =5802789;
#20;
$display("Result = %d", result); assert(result ==11864570);
row = 79;
ciphertext_entry =8048348;
#20;
$display("Result = %d", result); assert(result ==5451845);
row = 80;
ciphertext_entry =2613732;
#20;
$display("Result = %d", result); assert(result ==11717955);
row = 81;
ciphertext_entry =13810549;
#20;
$display("Result = %d", result); assert(result ==4129897);
row = 82;
ciphertext_entry =1025754;
#20;
$display("Result = %d", result); assert(result ==8149442);
row = 83;
ciphertext_entry =1300761;
#20;
$display("Result = %d", result); assert(result ==7141269);
row = 84;
ciphertext_entry =14396277;
#20;
$display("Result = %d", result); assert(result ==4339341);
row = 85;
ciphertext_entry =13247639;
#20;
$display("Result = %d", result); assert(result ==15181080);
row = 86;
ciphertext_entry =7378534;
#20;
$display("Result = %d", result); assert(result ==13676305);
row = 87;
ciphertext_entry =13578534;
#20;
$display("Result = %d", result); assert(result ==16333087);
row = 88;
ciphertext_entry =6631803;
#20;
$display("Result = %d", result); assert(result ==2421015);
row = 89;
ciphertext_entry =6539247;
#20;
$display("Result = %d", result); assert(result ==13393385);
row = 90;
ciphertext_entry =9670700;
#20;
$display("Result = %d", result); assert(result ==8002599);
row = 91;
ciphertext_entry =12541800;
#20;
$display("Result = %d", result); assert(result ==14313680);
row = 92;
ciphertext_entry =662742;
#20;
$display("Result = %d", result); assert(result ==2748062);
row = 93;
ciphertext_entry =14810215;
#20;
$display("Result = %d", result); assert(result ==10812337);
row = 94;
ciphertext_entry =14564306;
#20;
$display("Result = %d", result); assert(result ==7345114);
row = 95;
ciphertext_entry =15812604;
#20;
$display("Result = %d", result); assert(result ==14317782);
row = 96;
ciphertext_entry =878920;
#20;
$display("Result = %d", result); assert(result ==5634820);
row = 97;
ciphertext_entry =1179072;
#20;
$display("Result = %d", result); assert(result ==9237991);
row = 98;
ciphertext_entry =11098319;
#20;
$display("Result = %d", result); assert(result ==11250598);
row = 99;
ciphertext_entry =6504697;
#20;
$display("Result = %d", result); assert(result ==6299102);
row = 100;
ciphertext_entry =5157978;
#20;
$display("Result = %d", result); assert(result ==3495451);
row = 101;
ciphertext_entry =6349629;
#20;
$display("Result = %d", result); assert(result ==13159777);
row = 102;
ciphertext_entry =3513589;
#20;
$display("Result = %d", result); assert(result ==14399930);
row = 103;
ciphertext_entry =9104225;
#20;
$display("Result = %d", result); assert(result ==10433239);
row = 104;
ciphertext_entry =14514092;
#20;
$display("Result = %d", result); assert(result ==15568329);
row = 105;
ciphertext_entry =435730;
#20;
$display("Result = %d", result); assert(result ==2921027);
row = 106;
ciphertext_entry =3124935;
#20;
$display("Result = %d", result); assert(result ==9130627);
row = 107;
ciphertext_entry =7082632;
#20;
$display("Result = %d", result); assert(result ==10986881);
row = 108;
ciphertext_entry =15306750;
#20;
$display("Result = %d", result); assert(result ==12605471);
row = 109;
ciphertext_entry =10252241;
#20;
$display("Result = %d", result); assert(result ==678157);
row = 110;
ciphertext_entry =1517219;
#20;
$display("Result = %d", result); assert(result ==12092711);
row = 111;
ciphertext_entry =12865329;
#20;
$display("Result = %d", result); assert(result ==9962123);
row = 112;
ciphertext_entry =6884282;
#20;
$display("Result = %d", result); assert(result ==12061362);
row = 113;
ciphertext_entry =16527876;
#20;
$display("Result = %d", result); assert(result ==15987475);
row = 114;
ciphertext_entry =4831239;
#20;
$display("Result = %d", result); assert(result ==10046435);
row = 115;
ciphertext_entry =13777612;
#20;
$display("Result = %d", result); assert(result ==12755201);
row = 116;
ciphertext_entry =9520487;
#20;
$display("Result = %d", result); assert(result ==38038);
row = 117;
ciphertext_entry =1068946;
#20;
$display("Result = %d", result); assert(result ==9042483);
row = 118;
ciphertext_entry =1295344;
#20;
$display("Result = %d", result); assert(result ==14616324);
row = 119;
ciphertext_entry =14240044;
#20;
$display("Result = %d", result); assert(result ==2716062);
row = 120;
ciphertext_entry =11943159;
#20;
$display("Result = %d", result); assert(result ==2460887);
row = 121;
ciphertext_entry =8016467;
#20;
$display("Result = %d", result); assert(result ==9180482);
row = 122;
ciphertext_entry =9559681;
#20;
$display("Result = %d", result); assert(result ==16474798);
row = 123;
ciphertext_entry =3361994;
#20;
$display("Result = %d", result); assert(result ==9988796);
row = 124;
ciphertext_entry =3826283;
#20;
$display("Result = %d", result); assert(result ==1677474);
row = 125;
ciphertext_entry =16026884;
#20;
$display("Result = %d", result); assert(result ==657554);
row = 126;
ciphertext_entry =15484096;
#20;
$display("Result = %d", result); assert(result ==12306628);
row = 127;
ciphertext_entry =562818;
#20;
$display("Result = %d", result); assert(result ==4339472);
row = 128;
ciphertext_entry =13170074;
#20;
$display("Result = %d", result); assert(result ==8531164);
ciphertext_select = 0;
row = 129;
#20;
$display("Result = %d", result); assert(result ==14358092);
row = 130;
#20;
$display("Result = %d", result); assert(result ==14462444);
row = 131;
#20;
$display("Result = %d", result); assert(result ==1951020);
row = 132;
#20;
$display("Result = %d", result); assert(result ==14016486);
row = 133;
#20;
$display("Result = %d", result); assert(result ==909498);
row = 134;
#20;
$display("Result = %d", result); assert(result ==14367649);
row = 135;
#20;
$display("Result = %d", result); assert(result ==7564939);
row = 136;
#20;
$display("Result = %d", result); assert(result ==16708636);
row = 137;
#20;
$display("Result = %d", result); assert(result ==367906);
row = 138;
#20;
$display("Result = %d", result); assert(result ==8145650);
row = 139;
#20;
$display("Result = %d", result); assert(result ==13694240);
row = 140;
#20;
$display("Result = %d", result); assert(result ==6815570);
row = 141;
#20;
$display("Result = %d", result); assert(result ==4935084);
row = 142;
#20;
$display("Result = %d", result); assert(result ==12489520);
row = 143;
#20;
$display("Result = %d", result); assert(result ==10458574);
row = 144;
#20;
$display("Result = %d", result); assert(result ==2340302);
row = 145;
#20;
$display("Result = %d", result); assert(result ==2232016);
row = 146;
#20;
$display("Result = %d", result); assert(result ==5288771);
row = 147;
#20;
$display("Result = %d", result); assert(result ==10980763);
row = 148;
#20;
$display("Result = %d", result); assert(result ==15853890);
row = 149;
#20;
$display("Result = %d", result); assert(result ==16132527);
row = 150;
#20;
$display("Result = %d", result); assert(result ==4787910);
row = 151;
#20;
$display("Result = %d", result); assert(result ==13373842);
row = 152;
#20;
$display("Result = %d", result); assert(result ==14822416);
row = 153;
#20;
$display("Result = %d", result); assert(result ==6817805);
row = 154;
#20;
$display("Result = %d", result); assert(result ==12942883);
row = 155;
#20;
$display("Result = %d", result); assert(result ==15942004);
row = 156;
#20;
$display("Result = %d", result); assert(result ==8758360);
row = 157;
#20;
$display("Result = %d", result); assert(result ==5295643);
row = 158;
#20;
$display("Result = %d", result); assert(result ==760592);
row = 159;
#20;
$display("Result = %d", result); assert(result ==8889156);
row = 160;
#20;
$display("Result = %d", result); assert(result ==66581);
row = 161;
#20;
$display("Result = %d", result); assert(result ==3791407);
row = 162;
#20;
$display("Result = %d", result); assert(result ==7259792);
row = 163;
#20;
$display("Result = %d", result); assert(result ==11302337);
row = 164;
#20;
$display("Result = %d", result); assert(result ==1914236);
row = 165;
#20;
$display("Result = %d", result); assert(result ==13877243);
row = 166;
#20;
$display("Result = %d", result); assert(result ==13765392);
row = 167;
#20;
$display("Result = %d", result); assert(result ==3179701);
row = 168;
#20;
$display("Result = %d", result); assert(result ==2442324);
row = 169;
#20;
$display("Result = %d", result); assert(result ==12866732);
row = 170;
#20;
$display("Result = %d", result); assert(result ==15567379);
row = 171;
#20;
$display("Result = %d", result); assert(result ==10958773);
row = 172;
#20;
$display("Result = %d", result); assert(result ==7799290);
row = 173;
#20;
$display("Result = %d", result); assert(result ==4020506);
row = 174;
#20;
$display("Result = %d", result); assert(result ==6581360);
row = 175;
#20;
$display("Result = %d", result); assert(result ==98501);
row = 176;
#20;
$display("Result = %d", result); assert(result ==2601292);
row = 177;
#20;
$display("Result = %d", result); assert(result ==9965920);
row = 178;
#20;
$display("Result = %d", result); assert(result ==9195985);
row = 179;
#20;
$display("Result = %d", result); assert(result ==10368014);
row = 180;
#20;
$display("Result = %d", result); assert(result ==12651246);
row = 181;
#20;
$display("Result = %d", result); assert(result ==3139764);
row = 182;
#20;
$display("Result = %d", result); assert(result ==11006474);
row = 183;
#20;
$display("Result = %d", result); assert(result ==4412718);
row = 184;
#20;
$display("Result = %d", result); assert(result ==16487574);
row = 185;
#20;
$display("Result = %d", result); assert(result ==133985);
row = 186;
#20;
$display("Result = %d", result); assert(result ==11699478);
row = 187;
#20;
$display("Result = %d", result); assert(result ==14404876);
row = 188;
#20;
$display("Result = %d", result); assert(result ==1889198);
row = 189;
#20;
$display("Result = %d", result); assert(result ==10043132);
row = 190;
#20;
$display("Result = %d", result); assert(result ==15692938);
row = 191;
#20;
$display("Result = %d", result); assert(result ==5595491);
row = 192;
#20;
$display("Result = %d", result); assert(result ==4924678);
row = 193;
#20;
$display("Result = %d", result); assert(result ==11881539);
row = 194;
#20;
$display("Result = %d", result); assert(result ==14262027);
row = 195;
#20;
$display("Result = %d", result); assert(result ==12998256);
row = 196;
#20;
$display("Result = %d", result); assert(result ==1338779);
row = 197;
#20;
$display("Result = %d", result); assert(result ==13219471);
row = 198;
#20;
$display("Result = %d", result); assert(result ==4979893);
row = 199;
#20;
$display("Result = %d", result); assert(result ==15754346);
row = 200;
#20;
$display("Result = %d", result); assert(result ==5533285);
row = 201;
#20;
$display("Result = %d", result); assert(result ==12463183);
row = 202;
#20;
$display("Result = %d", result); assert(result ==15285131);
row = 203;
#20;
$display("Result = %d", result); assert(result ==12556576);
row = 204;
#20;
$display("Result = %d", result); assert(result ==15340824);
row = 205;
#20;
$display("Result = %d", result); assert(result ==8230660);
row = 206;
#20;
$display("Result = %d", result); assert(result ==10006947);
row = 207;
#20;
$display("Result = %d", result); assert(result ==6363531);
row = 208;
#20;
$display("Result = %d", result); assert(result ==16651766);
row = 209;
#20;
$display("Result = %d", result); assert(result ==1371245);
row = 210;
#20;
$display("Result = %d", result); assert(result ==14755683);
row = 211;
#20;
$display("Result = %d", result); assert(result ==40638);
row = 212;
#20;
$display("Result = %d", result); assert(result ==6770164);
row = 213;
#20;
$display("Result = %d", result); assert(result ==15713);
row = 214;
#20;
$display("Result = %d", result); assert(result ==5522971);
row = 215;
#20;
$display("Result = %d", result); assert(result ==879140);
row = 216;
#20;
$display("Result = %d", result); assert(result ==13973131);
row = 217;
#20;
$display("Result = %d", result); assert(result ==13465729);
row = 218;
#20;
$display("Result = %d", result); assert(result ==15017507);
row = 219;
#20;
$display("Result = %d", result); assert(result ==8032671);
row = 220;
#20;
$display("Result = %d", result); assert(result ==10029070);
row = 221;
#20;
$display("Result = %d", result); assert(result ==15128655);
row = 222;
#20;
$display("Result = %d", result); assert(result ==637274);
row = 223;
#20;
$display("Result = %d", result); assert(result ==9714436);
row = 224;
#20;
$display("Result = %d", result); assert(result ==1592235);
row = 225;
#20;
$display("Result = %d", result); assert(result ==16600251);
row = 226;
#20;
$display("Result = %d", result); assert(result ==12607184);
row = 227;
#20;
$display("Result = %d", result); assert(result ==1645089);
row = 228;
#20;
$display("Result = %d", result); assert(result ==16671604);
row = 229;
#20;
$display("Result = %d", result); assert(result ==3415124);
row = 230;
#20;
$display("Result = %d", result); assert(result ==1568361);
row = 231;
#20;
$display("Result = %d", result); assert(result ==1646623);
row = 232;
#20;
$display("Result = %d", result); assert(result ==9285577);
row = 233;
#20;
$display("Result = %d", result); assert(result ==6745648);
row = 234;
#20;
$display("Result = %d", result); assert(result ==14289563);
row = 235;
#20;
$display("Result = %d", result); assert(result ==14355712);
row = 236;
#20;
$display("Result = %d", result); assert(result ==919244);
row = 237;
#20;
$display("Result = %d", result); assert(result ==14982079);
row = 238;
#20;
$display("Result = %d", result); assert(result ==5961354);
row = 239;
#20;
$display("Result = %d", result); assert(result ==15270253);
row = 240;
#20;
$display("Result = %d", result); assert(result ==4528588);
row = 241;
#20;
$display("Result = %d", result); assert(result ==6033654);
row = 242;
#20;
$display("Result = %d", result); assert(result ==16753955);
row = 243;
#20;
$display("Result = %d", result); assert(result ==10808819);
row = 244;
#20;
$display("Result = %d", result); assert(result ==8803769);
row = 245;
#20;
$display("Result = %d", result); assert(result ==12401959);
row = 246;
#20;
$display("Result = %d", result); assert(result ==11366528);
row = 247;
#20;
$display("Result = %d", result); assert(result ==16490749);
row = 248;
#20;
$display("Result = %d", result); assert(result ==1561443);
row = 249;
#20;
$display("Result = %d", result); assert(result ==9690896);
row = 250;
#20;
$display("Result = %d", result); assert(result ==7419887);
row = 251;
#20;
$display("Result = %d", result); assert(result ==8895521);
row = 252;
#20;
$display("Result = %d", result); assert(result ==11099778);
row = 253;
#20;
$display("Result = %d", result); assert(result ==1480960);
row = 254;
#20;
$display("Result = %d", result); assert(result ==820600);
row = 255;
#20;
$display("Result = %d", result); assert(result ==16034846);
row = 256;
#20;
$display("Result = %d", result); assert(result ==16310052);
en=0;
rst_n=0;
#100;
rst_n=1;
#100;
en=1;
#20;
ciphertext_select = 0;
row = 0;
ciphertext_entry =5211550;
#20;
row = 1;
ciphertext_entry =14688493;
#20;
row = 2;
ciphertext_entry =13515507;
#20;
row = 3;
ciphertext_entry =10223486;
#20;
row = 4;
ciphertext_entry =15948488;
#20;
row = 5;
ciphertext_entry =15241648;
#20;
row = 6;
ciphertext_entry =6500362;
#20;
row = 7;
ciphertext_entry =4886935;
#20;
row = 8;
ciphertext_entry =13140336;
#20;
row = 9;
ciphertext_entry =8387096;
#20;
row = 10;
ciphertext_entry =16498127;
#20;
row = 11;
ciphertext_entry =15301879;
#20;
row = 12;
ciphertext_entry =1049822;
#20;
row = 13;
ciphertext_entry =16247570;
#20;
row = 14;
ciphertext_entry =175255;
#20;
row = 15;
ciphertext_entry =7862548;
#20;
row = 16;
ciphertext_entry =15783823;
#20;
row = 17;
ciphertext_entry =5740321;
#20;
row = 18;
ciphertext_entry =15284067;
#20;
row = 19;
ciphertext_entry =3862071;
#20;
row = 20;
ciphertext_entry =11986665;
#20;
row = 21;
ciphertext_entry =6820803;
#20;
row = 22;
ciphertext_entry =1904184;
#20;
row = 23;
ciphertext_entry =2497663;
#20;
row = 24;
ciphertext_entry =6474940;
#20;
row = 25;
ciphertext_entry =10468088;
#20;
row = 26;
ciphertext_entry =1184098;
#20;
row = 27;
ciphertext_entry =11560700;
#20;
row = 28;
ciphertext_entry =1749491;
#20;
row = 29;
ciphertext_entry =8495382;
#20;
row = 30;
ciphertext_entry =15909629;
#20;
row = 31;
ciphertext_entry =9693910;
#20;
row = 32;
ciphertext_entry =1239378;
#20;
row = 33;
ciphertext_entry =9024400;
#20;
row = 34;
ciphertext_entry =38293;
#20;
row = 35;
ciphertext_entry =15177299;
#20;
row = 36;
ciphertext_entry =15731280;
#20;
row = 37;
ciphertext_entry =13001685;
#20;
row = 38;
ciphertext_entry =542439;
#20;
row = 39;
ciphertext_entry =10524192;
#20;
row = 40;
ciphertext_entry =2291556;
#20;
row = 41;
ciphertext_entry =12408703;
#20;
row = 42;
ciphertext_entry =4190037;
#20;
row = 43;
ciphertext_entry =12734289;
#20;
row = 44;
ciphertext_entry =6001520;
#20;
row = 45;
ciphertext_entry =9137878;
#20;
row = 46;
ciphertext_entry =12664790;
#20;
row = 47;
ciphertext_entry =7124776;
#20;
row = 48;
ciphertext_entry =10140883;
#20;
row = 49;
ciphertext_entry =1270124;
#20;
row = 50;
ciphertext_entry =7214171;
#20;
row = 51;
ciphertext_entry =16211493;
#20;
row = 52;
ciphertext_entry =3708837;
#20;
row = 53;
ciphertext_entry =5259555;
#20;
row = 54;
ciphertext_entry =8313106;
#20;
row = 55;
ciphertext_entry =4578930;
#20;
row = 56;
ciphertext_entry =5152964;
#20;
row = 57;
ciphertext_entry =3398925;
#20;
row = 58;
ciphertext_entry =1172283;
#20;
row = 59;
ciphertext_entry =2998373;
#20;
row = 60;
ciphertext_entry =9376963;
#20;
row = 61;
ciphertext_entry =3865257;
#20;
row = 62;
ciphertext_entry =13693128;
#20;
row = 63;
ciphertext_entry =10592138;
#20;
row = 64;
ciphertext_entry =6115032;
#20;
row = 65;
ciphertext_entry =6527344;
#20;
row = 66;
ciphertext_entry =15565028;
#20;
row = 67;
ciphertext_entry =14395283;
#20;
row = 68;
ciphertext_entry =13113328;
#20;
row = 69;
ciphertext_entry =6788952;
#20;
row = 70;
ciphertext_entry =5808183;
#20;
row = 71;
ciphertext_entry =6643775;
#20;
row = 72;
ciphertext_entry =12126090;
#20;
row = 73;
ciphertext_entry =10264096;
#20;
row = 74;
ciphertext_entry =1020869;
#20;
row = 75;
ciphertext_entry =648941;
#20;
row = 76;
ciphertext_entry =14750184;
#20;
row = 77;
ciphertext_entry =12939364;
#20;
row = 78;
ciphertext_entry =12073190;
#20;
row = 79;
ciphertext_entry =16035452;
#20;
row = 80;
ciphertext_entry =15002556;
#20;
row = 81;
ciphertext_entry =15736732;
#20;
row = 82;
ciphertext_entry =4529541;
#20;
row = 83;
ciphertext_entry =11802161;
#20;
row = 84;
ciphertext_entry =2553561;
#20;
row = 85;
ciphertext_entry =5123961;
#20;
row = 86;
ciphertext_entry =8592169;
#20;
row = 87;
ciphertext_entry =2250872;
#20;
row = 88;
ciphertext_entry =656029;
#20;
row = 89;
ciphertext_entry =742801;
#20;
row = 90;
ciphertext_entry =729570;
#20;
row = 91;
ciphertext_entry =14916029;
#20;
row = 92;
ciphertext_entry =5210822;
#20;
row = 93;
ciphertext_entry =16411051;
#20;
row = 94;
ciphertext_entry =9019593;
#20;
row = 95;
ciphertext_entry =10693092;
#20;
row = 96;
ciphertext_entry =6304794;
#20;
row = 97;
ciphertext_entry =11521193;
#20;
row = 98;
ciphertext_entry =9032572;
#20;
row = 99;
ciphertext_entry =13387627;
#20;
row = 100;
ciphertext_entry =3263700;
#20;
row = 101;
ciphertext_entry =14937233;
#20;
row = 102;
ciphertext_entry =7429110;
#20;
row = 103;
ciphertext_entry =13232035;
#20;
row = 104;
ciphertext_entry =14859307;
#20;
row = 105;
ciphertext_entry =5602419;
#20;
row = 106;
ciphertext_entry =5306147;
#20;
row = 107;
ciphertext_entry =266145;
#20;
row = 108;
ciphertext_entry =5830760;
#20;
row = 109;
ciphertext_entry =16636288;
#20;
row = 110;
ciphertext_entry =1435555;
#20;
row = 111;
ciphertext_entry =14348898;
#20;
row = 112;
ciphertext_entry =13259936;
#20;
row = 113;
ciphertext_entry =2575570;
#20;
row = 114;
ciphertext_entry =15605249;
#20;
row = 115;
ciphertext_entry =4937508;
#20;
row = 116;
ciphertext_entry =9369569;
#20;
row = 117;
ciphertext_entry =1562993;
#20;
row = 118;
ciphertext_entry =15310888;
#20;
row = 119;
ciphertext_entry =498492;
#20;
row = 120;
ciphertext_entry =10919398;
#20;
row = 121;
ciphertext_entry =4919097;
#20;
row = 122;
ciphertext_entry =6840257;
#20;
row = 123;
ciphertext_entry =8048857;
#20;
row = 124;
ciphertext_entry =122956;
#20;
row = 125;
ciphertext_entry =5670519;
#20;
row = 126;
ciphertext_entry =6420922;
#20;
row = 127;
ciphertext_entry =7560556;
#20;
row = 128;
ciphertext_entry =532636;
#20;
ciphertext_select = 1;
row = 0;
ciphertext_entry =5211550;
#20;
$display("Result = %d", result); assert(result ==8712906);
row = 1;
ciphertext_entry =14688493;
#20;
$display("Result = %d", result); assert(result ==1973635);
row = 2;
ciphertext_entry =13515507;
#20;
$display("Result = %d", result); assert(result ==149851);
row = 3;
ciphertext_entry =10223486;
#20;
$display("Result = %d", result); assert(result ==13512620);
row = 4;
ciphertext_entry =15948488;
#20;
$display("Result = %d", result); assert(result ==14975511);
row = 5;
ciphertext_entry =15241648;
#20;
$display("Result = %d", result); assert(result ==10994961);
row = 6;
ciphertext_entry =6500362;
#20;
$display("Result = %d", result); assert(result ==4988679);
row = 7;
ciphertext_entry =4886935;
#20;
$display("Result = %d", result); assert(result ==3783264);
row = 8;
ciphertext_entry =13140336;
#20;
$display("Result = %d", result); assert(result ==10617830);
row = 9;
ciphertext_entry =8387096;
#20;
$display("Result = %d", result); assert(result ==15643446);
row = 10;
ciphertext_entry =16498127;
#20;
$display("Result = %d", result); assert(result ==16589587);
row = 11;
ciphertext_entry =15301879;
#20;
$display("Result = %d", result); assert(result ==3920008);
row = 12;
ciphertext_entry =1049822;
#20;
$display("Result = %d", result); assert(result ==8944932);
row = 13;
ciphertext_entry =16247570;
#20;
$display("Result = %d", result); assert(result ==11088622);
row = 14;
ciphertext_entry =175255;
#20;
$display("Result = %d", result); assert(result ==7209733);
row = 15;
ciphertext_entry =7862548;
#20;
$display("Result = %d", result); assert(result ==4465315);
row = 16;
ciphertext_entry =15783823;
#20;
$display("Result = %d", result); assert(result ==14946755);
row = 17;
ciphertext_entry =5740321;
#20;
$display("Result = %d", result); assert(result ==14206054);
row = 18;
ciphertext_entry =15284067;
#20;
$display("Result = %d", result); assert(result ==332220);
row = 19;
ciphertext_entry =3862071;
#20;
$display("Result = %d", result); assert(result ==10520310);
row = 20;
ciphertext_entry =11986665;
#20;
$display("Result = %d", result); assert(result ==7198140);
row = 21;
ciphertext_entry =6820803;
#20;
$display("Result = %d", result); assert(result ==10784301);
row = 22;
ciphertext_entry =1904184;
#20;
$display("Result = %d", result); assert(result ==3809779);
row = 23;
ciphertext_entry =2497663;
#20;
$display("Result = %d", result); assert(result ==15989273);
row = 24;
ciphertext_entry =6474940;
#20;
$display("Result = %d", result); assert(result ==1045977);
row = 25;
ciphertext_entry =10468088;
#20;
$display("Result = %d", result); assert(result ==12627093);
row = 26;
ciphertext_entry =1184098;
#20;
$display("Result = %d", result); assert(result ==9951190);
row = 27;
ciphertext_entry =11560700;
#20;
$display("Result = %d", result); assert(result ==6270535);
row = 28;
ciphertext_entry =1749491;
#20;
$display("Result = %d", result); assert(result ==14882761);
row = 29;
ciphertext_entry =8495382;
#20;
$display("Result = %d", result); assert(result ==5157090);
row = 30;
ciphertext_entry =15909629;
#20;
$display("Result = %d", result); assert(result ==7778953);
row = 31;
ciphertext_entry =9693910;
#20;
$display("Result = %d", result); assert(result ==10913963);
row = 32;
ciphertext_entry =1239378;
#20;
$display("Result = %d", result); assert(result ==15422453);
row = 33;
ciphertext_entry =9024400;
#20;
$display("Result = %d", result); assert(result ==6293765);
row = 34;
ciphertext_entry =38293;
#20;
$display("Result = %d", result); assert(result ==13035127);
row = 35;
ciphertext_entry =15177299;
#20;
$display("Result = %d", result); assert(result ==16501327);
row = 36;
ciphertext_entry =15731280;
#20;
$display("Result = %d", result); assert(result ==14765971);
row = 37;
ciphertext_entry =13001685;
#20;
$display("Result = %d", result); assert(result ==14493392);
row = 38;
ciphertext_entry =542439;
#20;
$display("Result = %d", result); assert(result ==10334508);
row = 39;
ciphertext_entry =10524192;
#20;
$display("Result = %d", result); assert(result ==12840221);
row = 40;
ciphertext_entry =2291556;
#20;
$display("Result = %d", result); assert(result ==10925059);
row = 41;
ciphertext_entry =12408703;
#20;
$display("Result = %d", result); assert(result ==811723);
row = 42;
ciphertext_entry =4190037;
#20;
$display("Result = %d", result); assert(result ==7368908);
row = 43;
ciphertext_entry =12734289;
#20;
$display("Result = %d", result); assert(result ==9265689);
row = 44;
ciphertext_entry =6001520;
#20;
$display("Result = %d", result); assert(result ==7569512);
row = 45;
ciphertext_entry =9137878;
#20;
$display("Result = %d", result); assert(result ==6644094);
row = 46;
ciphertext_entry =12664790;
#20;
$display("Result = %d", result); assert(result ==1613401);
row = 47;
ciphertext_entry =7124776;
#20;
$display("Result = %d", result); assert(result ==3544995);
row = 48;
ciphertext_entry =10140883;
#20;
$display("Result = %d", result); assert(result ==7705195);
row = 49;
ciphertext_entry =1270124;
#20;
$display("Result = %d", result); assert(result ==16140989);
row = 50;
ciphertext_entry =7214171;
#20;
$display("Result = %d", result); assert(result ==13419532);
row = 51;
ciphertext_entry =16211493;
#20;
$display("Result = %d", result); assert(result ==4634535);
row = 52;
ciphertext_entry =3708837;
#20;
$display("Result = %d", result); assert(result ==3452834);
row = 53;
ciphertext_entry =5259555;
#20;
$display("Result = %d", result); assert(result ==15683146);
row = 54;
ciphertext_entry =8313106;
#20;
$display("Result = %d", result); assert(result ==105106);
row = 55;
ciphertext_entry =4578930;
#20;
$display("Result = %d", result); assert(result ==7331326);
row = 56;
ciphertext_entry =5152964;
#20;
$display("Result = %d", result); assert(result ==4101226);
row = 57;
ciphertext_entry =3398925;
#20;
$display("Result = %d", result); assert(result ==13102277);
row = 58;
ciphertext_entry =1172283;
#20;
$display("Result = %d", result); assert(result ==12110923);
row = 59;
ciphertext_entry =2998373;
#20;
$display("Result = %d", result); assert(result ==14461994);
row = 60;
ciphertext_entry =9376963;
#20;
$display("Result = %d", result); assert(result ==7280429);
row = 61;
ciphertext_entry =3865257;
#20;
$display("Result = %d", result); assert(result ==8165063);
row = 62;
ciphertext_entry =13693128;
#20;
$display("Result = %d", result); assert(result ==779882);
row = 63;
ciphertext_entry =10592138;
#20;
$display("Result = %d", result); assert(result ==11728255);
row = 64;
ciphertext_entry =6115032;
#20;
$display("Result = %d", result); assert(result ==6337580);
row = 65;
ciphertext_entry =6527344;
#20;
$display("Result = %d", result); assert(result ==2032771);
row = 66;
ciphertext_entry =15565028;
#20;
$display("Result = %d", result); assert(result ==5171066);
row = 67;
ciphertext_entry =14395283;
#20;
$display("Result = %d", result); assert(result ==11425803);
row = 68;
ciphertext_entry =13113328;
#20;
$display("Result = %d", result); assert(result ==1276656);
row = 69;
ciphertext_entry =6788952;
#20;
$display("Result = %d", result); assert(result ==7963740);
row = 70;
ciphertext_entry =5808183;
#20;
$display("Result = %d", result); assert(result ==4915744);
row = 71;
ciphertext_entry =6643775;
#20;
$display("Result = %d", result); assert(result ==12078470);
row = 72;
ciphertext_entry =12126090;
#20;
$display("Result = %d", result); assert(result ==2265099);
row = 73;
ciphertext_entry =10264096;
#20;
$display("Result = %d", result); assert(result ==598974);
row = 74;
ciphertext_entry =1020869;
#20;
$display("Result = %d", result); assert(result ==14173803);
row = 75;
ciphertext_entry =648941;
#20;
$display("Result = %d", result); assert(result ==7955637);
row = 76;
ciphertext_entry =14750184;
#20;
$display("Result = %d", result); assert(result ==13479950);
row = 77;
ciphertext_entry =12939364;
#20;
$display("Result = %d", result); assert(result ==6698512);
row = 78;
ciphertext_entry =12073190;
#20;
$display("Result = %d", result); assert(result ==14068045);
row = 79;
ciphertext_entry =16035452;
#20;
$display("Result = %d", result); assert(result ==2373384);
row = 80;
ciphertext_entry =15002556;
#20;
$display("Result = %d", result); assert(result ==5629519);
row = 81;
ciphertext_entry =15736732;
#20;
$display("Result = %d", result); assert(result ==14492052);
row = 82;
ciphertext_entry =4529541;
#20;
$display("Result = %d", result); assert(result ==1679982);
row = 83;
ciphertext_entry =11802161;
#20;
$display("Result = %d", result); assert(result ==11348384);
row = 84;
ciphertext_entry =2553561;
#20;
$display("Result = %d", result); assert(result ==10924015);
row = 85;
ciphertext_entry =5123961;
#20;
$display("Result = %d", result); assert(result ==16134810);
row = 86;
ciphertext_entry =8592169;
#20;
$display("Result = %d", result); assert(result ==11318545);
row = 87;
ciphertext_entry =2250872;
#20;
$display("Result = %d", result); assert(result ==16448086);
row = 88;
ciphertext_entry =656029;
#20;
$display("Result = %d", result); assert(result ==9973341);
row = 89;
ciphertext_entry =742801;
#20;
$display("Result = %d", result); assert(result ==3204407);
row = 90;
ciphertext_entry =729570;
#20;
$display("Result = %d", result); assert(result ==10254961);
row = 91;
ciphertext_entry =14916029;
#20;
$display("Result = %d", result); assert(result ==14705348);
row = 92;
ciphertext_entry =5210822;
#20;
$display("Result = %d", result); assert(result ==4298260);
row = 93;
ciphertext_entry =16411051;
#20;
$display("Result = %d", result); assert(result ==2741539);
row = 94;
ciphertext_entry =9019593;
#20;
$display("Result = %d", result); assert(result ==1704230);
row = 95;
ciphertext_entry =10693092;
#20;
$display("Result = %d", result); assert(result ==9387937);
row = 96;
ciphertext_entry =6304794;
#20;
$display("Result = %d", result); assert(result ==2720992);
row = 97;
ciphertext_entry =11521193;
#20;
$display("Result = %d", result); assert(result ==11489309);
row = 98;
ciphertext_entry =9032572;
#20;
$display("Result = %d", result); assert(result ==16109135);
row = 99;
ciphertext_entry =13387627;
#20;
$display("Result = %d", result); assert(result ==6199972);
row = 100;
ciphertext_entry =3263700;
#20;
$display("Result = %d", result); assert(result ==7665882);
row = 101;
ciphertext_entry =14937233;
#20;
$display("Result = %d", result); assert(result ==16163228);
row = 102;
ciphertext_entry =7429110;
#20;
$display("Result = %d", result); assert(result ==909600);
row = 103;
ciphertext_entry =13232035;
#20;
$display("Result = %d", result); assert(result ==10586846);
row = 104;
ciphertext_entry =14859307;
#20;
$display("Result = %d", result); assert(result ==2561156);
row = 105;
ciphertext_entry =5602419;
#20;
$display("Result = %d", result); assert(result ==14980668);
row = 106;
ciphertext_entry =5306147;
#20;
$display("Result = %d", result); assert(result ==3698069);
row = 107;
ciphertext_entry =266145;
#20;
$display("Result = %d", result); assert(result ==16168960);
row = 108;
ciphertext_entry =5830760;
#20;
$display("Result = %d", result); assert(result ==10952380);
row = 109;
ciphertext_entry =16636288;
#20;
$display("Result = %d", result); assert(result ==1064579);
row = 110;
ciphertext_entry =1435555;
#20;
$display("Result = %d", result); assert(result ==15043526);
row = 111;
ciphertext_entry =14348898;
#20;
$display("Result = %d", result); assert(result ==458426);
row = 112;
ciphertext_entry =13259936;
#20;
$display("Result = %d", result); assert(result ==170649);
row = 113;
ciphertext_entry =2575570;
#20;
$display("Result = %d", result); assert(result ==14452801);
row = 114;
ciphertext_entry =15605249;
#20;
$display("Result = %d", result); assert(result ==12083960);
row = 115;
ciphertext_entry =4937508;
#20;
$display("Result = %d", result); assert(result ==6027319);
row = 116;
ciphertext_entry =9369569;
#20;
$display("Result = %d", result); assert(result ==15405321);
row = 117;
ciphertext_entry =1562993;
#20;
$display("Result = %d", result); assert(result ==14601939);
row = 118;
ciphertext_entry =15310888;
#20;
$display("Result = %d", result); assert(result ==11203383);
row = 119;
ciphertext_entry =498492;
#20;
$display("Result = %d", result); assert(result ==15507635);
row = 120;
ciphertext_entry =10919398;
#20;
$display("Result = %d", result); assert(result ==15303219);
row = 121;
ciphertext_entry =4919097;
#20;
$display("Result = %d", result); assert(result ==12410820);
row = 122;
ciphertext_entry =6840257;
#20;
$display("Result = %d", result); assert(result ==8065647);
row = 123;
ciphertext_entry =8048857;
#20;
$display("Result = %d", result); assert(result ==16750059);
row = 124;
ciphertext_entry =122956;
#20;
$display("Result = %d", result); assert(result ==693511);
row = 125;
ciphertext_entry =5670519;
#20;
$display("Result = %d", result); assert(result ==8819798);
row = 126;
ciphertext_entry =6420922;
#20;
$display("Result = %d", result); assert(result ==10565651);
row = 127;
ciphertext_entry =7560556;
#20;
$display("Result = %d", result); assert(result ==9997153);
row = 128;
ciphertext_entry =532636;
#20;
$display("Result = %d", result); assert(result ==8498519);
ciphertext_select = 0;
row = 129;
#20;
$display("Result = %d", result); assert(result ==5903063);
row = 130;
#20;
$display("Result = %d", result); assert(result ==3697251);
row = 131;
#20;
$display("Result = %d", result); assert(result ==16219931);
row = 132;
#20;
$display("Result = %d", result); assert(result ==11769545);
row = 133;
#20;
$display("Result = %d", result); assert(result ==10502036);
row = 134;
#20;
$display("Result = %d", result); assert(result ==12527066);
row = 135;
#20;
$display("Result = %d", result); assert(result ==14108806);
row = 136;
#20;
$display("Result = %d", result); assert(result ==14756257);
row = 137;
#20;
$display("Result = %d", result); assert(result ==8519341);
row = 138;
#20;
$display("Result = %d", result); assert(result ==2921207);
row = 139;
#20;
$display("Result = %d", result); assert(result ==1097574);
row = 140;
#20;
$display("Result = %d", result); assert(result ==5152114);
row = 141;
#20;
$display("Result = %d", result); assert(result ==4847763);
row = 142;
#20;
$display("Result = %d", result); assert(result ==9593228);
row = 143;
#20;
$display("Result = %d", result); assert(result ==12794040);
row = 144;
#20;
$display("Result = %d", result); assert(result ==15723466);
row = 145;
#20;
$display("Result = %d", result); assert(result ==7034334);
row = 146;
#20;
$display("Result = %d", result); assert(result ==5339051);
row = 147;
#20;
$display("Result = %d", result); assert(result ==8478389);
row = 148;
#20;
$display("Result = %d", result); assert(result ==11740721);
row = 149;
#20;
$display("Result = %d", result); assert(result ==815642);
row = 150;
#20;
$display("Result = %d", result); assert(result ==37126);
row = 151;
#20;
$display("Result = %d", result); assert(result ==9653586);
row = 152;
#20;
$display("Result = %d", result); assert(result ==5263854);
row = 153;
#20;
$display("Result = %d", result); assert(result ==16499383);
row = 154;
#20;
$display("Result = %d", result); assert(result ==4615820);
row = 155;
#20;
$display("Result = %d", result); assert(result ==9233368);
row = 156;
#20;
$display("Result = %d", result); assert(result ==11071180);
row = 157;
#20;
$display("Result = %d", result); assert(result ==6544624);
row = 158;
#20;
$display("Result = %d", result); assert(result ==7781661);
row = 159;
#20;
$display("Result = %d", result); assert(result ==4239380);
row = 160;
#20;
$display("Result = %d", result); assert(result ==6685728);
row = 161;
#20;
$display("Result = %d", result); assert(result ==12658378);
row = 162;
#20;
$display("Result = %d", result); assert(result ==5314895);
row = 163;
#20;
$display("Result = %d", result); assert(result ==9301633);
row = 164;
#20;
$display("Result = %d", result); assert(result ==4253661);
row = 165;
#20;
$display("Result = %d", result); assert(result ==10339381);
row = 166;
#20;
$display("Result = %d", result); assert(result ==1358067);
row = 167;
#20;
$display("Result = %d", result); assert(result ==2867938);
row = 168;
#20;
$display("Result = %d", result); assert(result ==14872994);
row = 169;
#20;
$display("Result = %d", result); assert(result ==11105826);
row = 170;
#20;
$display("Result = %d", result); assert(result ==2003035);
row = 171;
#20;
$display("Result = %d", result); assert(result ==2802571);
row = 172;
#20;
$display("Result = %d", result); assert(result ==11938573);
row = 173;
#20;
$display("Result = %d", result); assert(result ==4196796);
row = 174;
#20;
$display("Result = %d", result); assert(result ==9107959);
row = 175;
#20;
$display("Result = %d", result); assert(result ==6506498);
row = 176;
#20;
$display("Result = %d", result); assert(result ==11888433);
row = 177;
#20;
$display("Result = %d", result); assert(result ==14180724);
row = 178;
#20;
$display("Result = %d", result); assert(result ==1081072);
row = 179;
#20;
$display("Result = %d", result); assert(result ==13827568);
row = 180;
#20;
$display("Result = %d", result); assert(result ==9561116);
row = 181;
#20;
$display("Result = %d", result); assert(result ==4272528);
row = 182;
#20;
$display("Result = %d", result); assert(result ==4778383);
row = 183;
#20;
$display("Result = %d", result); assert(result ==11596203);
row = 184;
#20;
$display("Result = %d", result); assert(result ==12432794);
row = 185;
#20;
$display("Result = %d", result); assert(result ==11300134);
row = 186;
#20;
$display("Result = %d", result); assert(result ==15323416);
row = 187;
#20;
$display("Result = %d", result); assert(result ==11790118);
row = 188;
#20;
$display("Result = %d", result); assert(result ==5146909);
row = 189;
#20;
$display("Result = %d", result); assert(result ==16119801);
row = 190;
#20;
$display("Result = %d", result); assert(result ==1672500);
row = 191;
#20;
$display("Result = %d", result); assert(result ==964835);
row = 192;
#20;
$display("Result = %d", result); assert(result ==3268358);
row = 193;
#20;
$display("Result = %d", result); assert(result ==10683801);
row = 194;
#20;
$display("Result = %d", result); assert(result ==10664827);
row = 195;
#20;
$display("Result = %d", result); assert(result ==16371582);
row = 196;
#20;
$display("Result = %d", result); assert(result ==14508774);
row = 197;
#20;
$display("Result = %d", result); assert(result ==16346868);
row = 198;
#20;
$display("Result = %d", result); assert(result ==8054043);
row = 199;
#20;
$display("Result = %d", result); assert(result ==13762886);
row = 200;
#20;
$display("Result = %d", result); assert(result ==13692484);
row = 201;
#20;
$display("Result = %d", result); assert(result ==7654459);
row = 202;
#20;
$display("Result = %d", result); assert(result ==9820919);
row = 203;
#20;
$display("Result = %d", result); assert(result ==8014933);
row = 204;
#20;
$display("Result = %d", result); assert(result ==14033597);
row = 205;
#20;
$display("Result = %d", result); assert(result ==15119183);
row = 206;
#20;
$display("Result = %d", result); assert(result ==8487922);
row = 207;
#20;
$display("Result = %d", result); assert(result ==8215658);
row = 208;
#20;
$display("Result = %d", result); assert(result ==5148826);
row = 209;
#20;
$display("Result = %d", result); assert(result ==3073088);
row = 210;
#20;
$display("Result = %d", result); assert(result ==8705149);
row = 211;
#20;
$display("Result = %d", result); assert(result ==11819613);
row = 212;
#20;
$display("Result = %d", result); assert(result ==14313358);
row = 213;
#20;
$display("Result = %d", result); assert(result ==7792984);
row = 214;
#20;
$display("Result = %d", result); assert(result ==10675526);
row = 215;
#20;
$display("Result = %d", result); assert(result ==4430275);
row = 216;
#20;
$display("Result = %d", result); assert(result ==12228682);
row = 217;
#20;
$display("Result = %d", result); assert(result ==16466173);
row = 218;
#20;
$display("Result = %d", result); assert(result ==9206901);
row = 219;
#20;
$display("Result = %d", result); assert(result ==15883979);
row = 220;
#20;
$display("Result = %d", result); assert(result ==14756566);
row = 221;
#20;
$display("Result = %d", result); assert(result ==14711089);
row = 222;
#20;
$display("Result = %d", result); assert(result ==15997232);
row = 223;
#20;
$display("Result = %d", result); assert(result ==457269);
row = 224;
#20;
$display("Result = %d", result); assert(result ==7968887);
row = 225;
#20;
$display("Result = %d", result); assert(result ==11468972);
row = 226;
#20;
$display("Result = %d", result); assert(result ==14326844);
row = 227;
#20;
$display("Result = %d", result); assert(result ==11173053);
row = 228;
#20;
$display("Result = %d", result); assert(result ==6058748);
row = 229;
#20;
$display("Result = %d", result); assert(result ==922718);
row = 230;
#20;
$display("Result = %d", result); assert(result ==7569439);
row = 231;
#20;
$display("Result = %d", result); assert(result ==6574531);
row = 232;
#20;
$display("Result = %d", result); assert(result ==5591825);
row = 233;
#20;
$display("Result = %d", result); assert(result ==2328714);
row = 234;
#20;
$display("Result = %d", result); assert(result ==7992875);
row = 235;
#20;
$display("Result = %d", result); assert(result ==4583585);
row = 236;
#20;
$display("Result = %d", result); assert(result ==11234521);
row = 237;
#20;
$display("Result = %d", result); assert(result ==12849125);
row = 238;
#20;
$display("Result = %d", result); assert(result ==3982359);
row = 239;
#20;
$display("Result = %d", result); assert(result ==11671016);
row = 240;
#20;
$display("Result = %d", result); assert(result ==14348097);
row = 241;
#20;
$display("Result = %d", result); assert(result ==7151660);
row = 242;
#20;
$display("Result = %d", result); assert(result ==1430175);
row = 243;
#20;
$display("Result = %d", result); assert(result ==6056267);
row = 244;
#20;
$display("Result = %d", result); assert(result ==2479057);
row = 245;
#20;
$display("Result = %d", result); assert(result ==12506101);
row = 246;
#20;
$display("Result = %d", result); assert(result ==1824843);
row = 247;
#20;
$display("Result = %d", result); assert(result ==10825531);
row = 248;
#20;
$display("Result = %d", result); assert(result ==11775852);
row = 249;
#20;
$display("Result = %d", result); assert(result ==11141919);
row = 250;
#20;
$display("Result = %d", result); assert(result ==15865467);
row = 251;
#20;
$display("Result = %d", result); assert(result ==12486464);
row = 252;
#20;
$display("Result = %d", result); assert(result ==5358702);
row = 253;
#20;
$display("Result = %d", result); assert(result ==14263966);
row = 254;
#20;
$display("Result = %d", result); assert(result ==3468444);
row = 255;
#20;
$display("Result = %d", result); assert(result ==16311280);
row = 256;
#20;
$display("Result = %d", result); assert(result ==16355736);
en=0;
rst_n=0;
#100;
rst_n=1;
#100;
en=1;
#20;
ciphertext_select = 0;
row = 0;
ciphertext_entry =10348332;
#20;
row = 1;
ciphertext_entry =16541935;
#20;
row = 2;
ciphertext_entry =6886586;
#20;
row = 3;
ciphertext_entry =2820101;
#20;
row = 4;
ciphertext_entry =12828906;
#20;
row = 5;
ciphertext_entry =10246417;
#20;
row = 6;
ciphertext_entry =5342173;
#20;
row = 7;
ciphertext_entry =11103339;
#20;
row = 8;
ciphertext_entry =6415174;
#20;
row = 9;
ciphertext_entry =15699522;
#20;
row = 10;
ciphertext_entry =1496028;
#20;
row = 11;
ciphertext_entry =13006037;
#20;
row = 12;
ciphertext_entry =16519691;
#20;
row = 13;
ciphertext_entry =7873607;
#20;
row = 14;
ciphertext_entry =10903096;
#20;
row = 15;
ciphertext_entry =10008768;
#20;
row = 16;
ciphertext_entry =9119507;
#20;
row = 17;
ciphertext_entry =10516517;
#20;
row = 18;
ciphertext_entry =14525461;
#20;
row = 19;
ciphertext_entry =4592326;
#20;
row = 20;
ciphertext_entry =15682335;
#20;
row = 21;
ciphertext_entry =3697395;
#20;
row = 22;
ciphertext_entry =13836424;
#20;
row = 23;
ciphertext_entry =3316229;
#20;
row = 24;
ciphertext_entry =10477501;
#20;
row = 25;
ciphertext_entry =7937268;
#20;
row = 26;
ciphertext_entry =1608395;
#20;
row = 27;
ciphertext_entry =15121414;
#20;
row = 28;
ciphertext_entry =1408979;
#20;
row = 29;
ciphertext_entry =231686;
#20;
row = 30;
ciphertext_entry =3906383;
#20;
row = 31;
ciphertext_entry =14744602;
#20;
row = 32;
ciphertext_entry =2515608;
#20;
row = 33;
ciphertext_entry =14090613;
#20;
row = 34;
ciphertext_entry =7164917;
#20;
row = 35;
ciphertext_entry =9337568;
#20;
row = 36;
ciphertext_entry =1884500;
#20;
row = 37;
ciphertext_entry =10266535;
#20;
row = 38;
ciphertext_entry =2628939;
#20;
row = 39;
ciphertext_entry =14376850;
#20;
row = 40;
ciphertext_entry =5708179;
#20;
row = 41;
ciphertext_entry =15444494;
#20;
row = 42;
ciphertext_entry =10383265;
#20;
row = 43;
ciphertext_entry =6552963;
#20;
row = 44;
ciphertext_entry =12614494;
#20;
row = 45;
ciphertext_entry =16428692;
#20;
row = 46;
ciphertext_entry =14536402;
#20;
row = 47;
ciphertext_entry =8807551;
#20;
row = 48;
ciphertext_entry =6016857;
#20;
row = 49;
ciphertext_entry =15880850;
#20;
row = 50;
ciphertext_entry =1437397;
#20;
row = 51;
ciphertext_entry =555166;
#20;
row = 52;
ciphertext_entry =6129311;
#20;
row = 53;
ciphertext_entry =3920652;
#20;
row = 54;
ciphertext_entry =2122950;
#20;
row = 55;
ciphertext_entry =4355986;
#20;
row = 56;
ciphertext_entry =13014627;
#20;
row = 57;
ciphertext_entry =8397752;
#20;
row = 58;
ciphertext_entry =12751183;
#20;
row = 59;
ciphertext_entry =1777770;
#20;
row = 60;
ciphertext_entry =10594057;
#20;
row = 61;
ciphertext_entry =15335468;
#20;
row = 62;
ciphertext_entry =1164330;
#20;
row = 63;
ciphertext_entry =7725848;
#20;
row = 64;
ciphertext_entry =6642888;
#20;
row = 65;
ciphertext_entry =6934284;
#20;
row = 66;
ciphertext_entry =3423927;
#20;
row = 67;
ciphertext_entry =2992075;
#20;
row = 68;
ciphertext_entry =10635199;
#20;
row = 69;
ciphertext_entry =3373210;
#20;
row = 70;
ciphertext_entry =1669468;
#20;
row = 71;
ciphertext_entry =4526647;
#20;
row = 72;
ciphertext_entry =12023394;
#20;
row = 73;
ciphertext_entry =2502984;
#20;
row = 74;
ciphertext_entry =11671049;
#20;
row = 75;
ciphertext_entry =15762439;
#20;
row = 76;
ciphertext_entry =15337319;
#20;
row = 77;
ciphertext_entry =6712255;
#20;
row = 78;
ciphertext_entry =631689;
#20;
row = 79;
ciphertext_entry =13104297;
#20;
row = 80;
ciphertext_entry =11043315;
#20;
row = 81;
ciphertext_entry =4371225;
#20;
row = 82;
ciphertext_entry =15753112;
#20;
row = 83;
ciphertext_entry =13422210;
#20;
row = 84;
ciphertext_entry =3353968;
#20;
row = 85;
ciphertext_entry =7849071;
#20;
row = 86;
ciphertext_entry =11929205;
#20;
row = 87;
ciphertext_entry =16329007;
#20;
row = 88;
ciphertext_entry =13086578;
#20;
row = 89;
ciphertext_entry =5710956;
#20;
row = 90;
ciphertext_entry =1862750;
#20;
row = 91;
ciphertext_entry =3848235;
#20;
row = 92;
ciphertext_entry =10222683;
#20;
row = 93;
ciphertext_entry =6359684;
#20;
row = 94;
ciphertext_entry =5148762;
#20;
row = 95;
ciphertext_entry =8900719;
#20;
row = 96;
ciphertext_entry =179002;
#20;
row = 97;
ciphertext_entry =394010;
#20;
row = 98;
ciphertext_entry =3835151;
#20;
row = 99;
ciphertext_entry =9792619;
#20;
row = 100;
ciphertext_entry =15930568;
#20;
row = 101;
ciphertext_entry =5758030;
#20;
row = 102;
ciphertext_entry =15213246;
#20;
row = 103;
ciphertext_entry =1110920;
#20;
row = 104;
ciphertext_entry =16043997;
#20;
row = 105;
ciphertext_entry =13051848;
#20;
row = 106;
ciphertext_entry =4867960;
#20;
row = 107;
ciphertext_entry =16168891;
#20;
row = 108;
ciphertext_entry =11594356;
#20;
row = 109;
ciphertext_entry =14898749;
#20;
row = 110;
ciphertext_entry =16349839;
#20;
row = 111;
ciphertext_entry =9019766;
#20;
row = 112;
ciphertext_entry =1249564;
#20;
row = 113;
ciphertext_entry =4337790;
#20;
row = 114;
ciphertext_entry =5514846;
#20;
row = 115;
ciphertext_entry =3026824;
#20;
row = 116;
ciphertext_entry =8097162;
#20;
row = 117;
ciphertext_entry =254588;
#20;
row = 118;
ciphertext_entry =13211275;
#20;
row = 119;
ciphertext_entry =5776563;
#20;
row = 120;
ciphertext_entry =2293504;
#20;
row = 121;
ciphertext_entry =11126760;
#20;
row = 122;
ciphertext_entry =2312572;
#20;
row = 123;
ciphertext_entry =16016002;
#20;
row = 124;
ciphertext_entry =12841246;
#20;
row = 125;
ciphertext_entry =7390091;
#20;
row = 126;
ciphertext_entry =16599182;
#20;
row = 127;
ciphertext_entry =16668189;
#20;
row = 128;
ciphertext_entry =1923577;
#20;
ciphertext_select = 1;
row = 0;
ciphertext_entry =10348332;
#20;
$display("Result = %d", result); assert(result ==13471776);
row = 1;
ciphertext_entry =16541935;
#20;
$display("Result = %d", result); assert(result ==16253088);
row = 2;
ciphertext_entry =6886586;
#20;
$display("Result = %d", result); assert(result ==10826142);
row = 3;
ciphertext_entry =2820101;
#20;
$display("Result = %d", result); assert(result ==8558742);
row = 4;
ciphertext_entry =12828906;
#20;
$display("Result = %d", result); assert(result ==10249611);
row = 5;
ciphertext_entry =10246417;
#20;
$display("Result = %d", result); assert(result ==1168603);
row = 6;
ciphertext_entry =5342173;
#20;
$display("Result = %d", result); assert(result ==14472918);
row = 7;
ciphertext_entry =11103339;
#20;
$display("Result = %d", result); assert(result ==16669532);
row = 8;
ciphertext_entry =6415174;
#20;
$display("Result = %d", result); assert(result ==12569082);
row = 9;
ciphertext_entry =15699522;
#20;
$display("Result = %d", result); assert(result ==6505524);
row = 10;
ciphertext_entry =1496028;
#20;
$display("Result = %d", result); assert(result ==9790746);
row = 11;
ciphertext_entry =13006037;
#20;
$display("Result = %d", result); assert(result ==12598684);
row = 12;
ciphertext_entry =16519691;
#20;
$display("Result = %d", result); assert(result ==9110911);
row = 13;
ciphertext_entry =7873607;
#20;
$display("Result = %d", result); assert(result ==8009683);
row = 14;
ciphertext_entry =10903096;
#20;
$display("Result = %d", result); assert(result ==16260914);
row = 15;
ciphertext_entry =10008768;
#20;
$display("Result = %d", result); assert(result ==16742215);
row = 16;
ciphertext_entry =9119507;
#20;
$display("Result = %d", result); assert(result ==6188902);
row = 17;
ciphertext_entry =10516517;
#20;
$display("Result = %d", result); assert(result ==8224417);
row = 18;
ciphertext_entry =14525461;
#20;
$display("Result = %d", result); assert(result ==11690500);
row = 19;
ciphertext_entry =4592326;
#20;
$display("Result = %d", result); assert(result ==411316);
row = 20;
ciphertext_entry =15682335;
#20;
$display("Result = %d", result); assert(result ==14928655);
row = 21;
ciphertext_entry =3697395;
#20;
$display("Result = %d", result); assert(result ==15035056);
row = 22;
ciphertext_entry =13836424;
#20;
$display("Result = %d", result); assert(result ==16211012);
row = 23;
ciphertext_entry =3316229;
#20;
$display("Result = %d", result); assert(result ==11114539);
row = 24;
ciphertext_entry =10477501;
#20;
$display("Result = %d", result); assert(result ==11106046);
row = 25;
ciphertext_entry =7937268;
#20;
$display("Result = %d", result); assert(result ==11812138);
row = 26;
ciphertext_entry =1608395;
#20;
$display("Result = %d", result); assert(result ==16282578);
row = 27;
ciphertext_entry =15121414;
#20;
$display("Result = %d", result); assert(result ==14094637);
row = 28;
ciphertext_entry =1408979;
#20;
$display("Result = %d", result); assert(result ==6345430);
row = 29;
ciphertext_entry =231686;
#20;
$display("Result = %d", result); assert(result ==16261000);
row = 30;
ciphertext_entry =3906383;
#20;
$display("Result = %d", result); assert(result ==8613451);
row = 31;
ciphertext_entry =14744602;
#20;
$display("Result = %d", result); assert(result ==1260808);
row = 32;
ciphertext_entry =2515608;
#20;
$display("Result = %d", result); assert(result ==1508190);
row = 33;
ciphertext_entry =14090613;
#20;
$display("Result = %d", result); assert(result ==9309113);
row = 34;
ciphertext_entry =7164917;
#20;
$display("Result = %d", result); assert(result ==13087282);
row = 35;
ciphertext_entry =9337568;
#20;
$display("Result = %d", result); assert(result ==9349889);
row = 36;
ciphertext_entry =1884500;
#20;
$display("Result = %d", result); assert(result ==6575375);
row = 37;
ciphertext_entry =10266535;
#20;
$display("Result = %d", result); assert(result ==12856079);
row = 38;
ciphertext_entry =2628939;
#20;
$display("Result = %d", result); assert(result ==975261);
row = 39;
ciphertext_entry =14376850;
#20;
$display("Result = %d", result); assert(result ==5298810);
row = 40;
ciphertext_entry =5708179;
#20;
$display("Result = %d", result); assert(result ==13921816);
row = 41;
ciphertext_entry =15444494;
#20;
$display("Result = %d", result); assert(result ==16737423);
row = 42;
ciphertext_entry =10383265;
#20;
$display("Result = %d", result); assert(result ==10917059);
row = 43;
ciphertext_entry =6552963;
#20;
$display("Result = %d", result); assert(result ==14944190);
row = 44;
ciphertext_entry =12614494;
#20;
$display("Result = %d", result); assert(result ==3027547);
row = 45;
ciphertext_entry =16428692;
#20;
$display("Result = %d", result); assert(result ==11231005);
row = 46;
ciphertext_entry =14536402;
#20;
$display("Result = %d", result); assert(result ==15250633);
row = 47;
ciphertext_entry =8807551;
#20;
$display("Result = %d", result); assert(result ==724809);
row = 48;
ciphertext_entry =6016857;
#20;
$display("Result = %d", result); assert(result ==2865431);
row = 49;
ciphertext_entry =15880850;
#20;
$display("Result = %d", result); assert(result ==16032657);
row = 50;
ciphertext_entry =1437397;
#20;
$display("Result = %d", result); assert(result ==7858762);
row = 51;
ciphertext_entry =555166;
#20;
$display("Result = %d", result); assert(result ==7725751);
row = 52;
ciphertext_entry =6129311;
#20;
$display("Result = %d", result); assert(result ==14181190);
row = 53;
ciphertext_entry =3920652;
#20;
$display("Result = %d", result); assert(result ==2174543);
row = 54;
ciphertext_entry =2122950;
#20;
$display("Result = %d", result); assert(result ==11734158);
row = 55;
ciphertext_entry =4355986;
#20;
$display("Result = %d", result); assert(result ==3054936);
row = 56;
ciphertext_entry =13014627;
#20;
$display("Result = %d", result); assert(result ==13431895);
row = 57;
ciphertext_entry =8397752;
#20;
$display("Result = %d", result); assert(result ==8961629);
row = 58;
ciphertext_entry =12751183;
#20;
$display("Result = %d", result); assert(result ==15610589);
row = 59;
ciphertext_entry =1777770;
#20;
$display("Result = %d", result); assert(result ==7146924);
row = 60;
ciphertext_entry =10594057;
#20;
$display("Result = %d", result); assert(result ==608882);
row = 61;
ciphertext_entry =15335468;
#20;
$display("Result = %d", result); assert(result ==8290717);
row = 62;
ciphertext_entry =1164330;
#20;
$display("Result = %d", result); assert(result ==13789829);
row = 63;
ciphertext_entry =7725848;
#20;
$display("Result = %d", result); assert(result ==15216086);
row = 64;
ciphertext_entry =6642888;
#20;
$display("Result = %d", result); assert(result ==8333858);
row = 65;
ciphertext_entry =6934284;
#20;
$display("Result = %d", result); assert(result ==8613557);
row = 66;
ciphertext_entry =3423927;
#20;
$display("Result = %d", result); assert(result ==10831700);
row = 67;
ciphertext_entry =2992075;
#20;
$display("Result = %d", result); assert(result ==5416556);
row = 68;
ciphertext_entry =10635199;
#20;
$display("Result = %d", result); assert(result ==3450490);
row = 69;
ciphertext_entry =3373210;
#20;
$display("Result = %d", result); assert(result ==15358844);
row = 70;
ciphertext_entry =1669468;
#20;
$display("Result = %d", result); assert(result ==16180472);
row = 71;
ciphertext_entry =4526647;
#20;
$display("Result = %d", result); assert(result ==7304623);
row = 72;
ciphertext_entry =12023394;
#20;
$display("Result = %d", result); assert(result ==15372758);
row = 73;
ciphertext_entry =2502984;
#20;
$display("Result = %d", result); assert(result ==9283588);
row = 74;
ciphertext_entry =11671049;
#20;
$display("Result = %d", result); assert(result ==922083);
row = 75;
ciphertext_entry =15762439;
#20;
$display("Result = %d", result); assert(result ==9966189);
row = 76;
ciphertext_entry =15337319;
#20;
$display("Result = %d", result); assert(result ==12548819);
row = 77;
ciphertext_entry =6712255;
#20;
$display("Result = %d", result); assert(result ==969413);
row = 78;
ciphertext_entry =631689;
#20;
$display("Result = %d", result); assert(result ==3217196);
row = 79;
ciphertext_entry =13104297;
#20;
$display("Result = %d", result); assert(result ==7664067);
row = 80;
ciphertext_entry =11043315;
#20;
$display("Result = %d", result); assert(result ==3353285);
row = 81;
ciphertext_entry =4371225;
#20;
$display("Result = %d", result); assert(result ==4658107);
row = 82;
ciphertext_entry =15753112;
#20;
$display("Result = %d", result); assert(result ==15133541);
row = 83;
ciphertext_entry =13422210;
#20;
$display("Result = %d", result); assert(result ==9578983);
row = 84;
ciphertext_entry =3353968;
#20;
$display("Result = %d", result); assert(result ==10249612);
row = 85;
ciphertext_entry =7849071;
#20;
$display("Result = %d", result); assert(result ==657228);
row = 86;
ciphertext_entry =11929205;
#20;
$display("Result = %d", result); assert(result ==1314898);
row = 87;
ciphertext_entry =16329007;
#20;
$display("Result = %d", result); assert(result ==11206009);
row = 88;
ciphertext_entry =13086578;
#20;
$display("Result = %d", result); assert(result ==3684410);
row = 89;
ciphertext_entry =5710956;
#20;
$display("Result = %d", result); assert(result ==16189694);
row = 90;
ciphertext_entry =1862750;
#20;
$display("Result = %d", result); assert(result ==5911906);
row = 91;
ciphertext_entry =3848235;
#20;
$display("Result = %d", result); assert(result ==1073607);
row = 92;
ciphertext_entry =10222683;
#20;
$display("Result = %d", result); assert(result ==12219197);
row = 93;
ciphertext_entry =6359684;
#20;
$display("Result = %d", result); assert(result ==7396039);
row = 94;
ciphertext_entry =5148762;
#20;
$display("Result = %d", result); assert(result ==12263636);
row = 95;
ciphertext_entry =8900719;
#20;
$display("Result = %d", result); assert(result ==14368716);
row = 96;
ciphertext_entry =179002;
#20;
$display("Result = %d", result); assert(result ==15458348);
row = 97;
ciphertext_entry =394010;
#20;
$display("Result = %d", result); assert(result ==8508379);
row = 98;
ciphertext_entry =3835151;
#20;
$display("Result = %d", result); assert(result ==12084478);
row = 99;
ciphertext_entry =9792619;
#20;
$display("Result = %d", result); assert(result ==15793090);
row = 100;
ciphertext_entry =15930568;
#20;
$display("Result = %d", result); assert(result ==1293800);
row = 101;
ciphertext_entry =5758030;
#20;
$display("Result = %d", result); assert(result ==12062577);
row = 102;
ciphertext_entry =15213246;
#20;
$display("Result = %d", result); assert(result ==2377676);
row = 103;
ciphertext_entry =1110920;
#20;
$display("Result = %d", result); assert(result ==212658);
row = 104;
ciphertext_entry =16043997;
#20;
$display("Result = %d", result); assert(result ==4855448);
row = 105;
ciphertext_entry =13051848;
#20;
$display("Result = %d", result); assert(result ==5823728);
row = 106;
ciphertext_entry =4867960;
#20;
$display("Result = %d", result); assert(result ==6828537);
row = 107;
ciphertext_entry =16168891;
#20;
$display("Result = %d", result); assert(result ==8999530);
row = 108;
ciphertext_entry =11594356;
#20;
$display("Result = %d", result); assert(result ==1181613);
row = 109;
ciphertext_entry =14898749;
#20;
$display("Result = %d", result); assert(result ==14690624);
row = 110;
ciphertext_entry =16349839;
#20;
$display("Result = %d", result); assert(result ==298795);
row = 111;
ciphertext_entry =9019766;
#20;
$display("Result = %d", result); assert(result ==1591336);
row = 112;
ciphertext_entry =1249564;
#20;
$display("Result = %d", result); assert(result ==13059748);
row = 113;
ciphertext_entry =4337790;
#20;
$display("Result = %d", result); assert(result ==12460786);
row = 114;
ciphertext_entry =5514846;
#20;
$display("Result = %d", result); assert(result ==5940592);
row = 115;
ciphertext_entry =3026824;
#20;
$display("Result = %d", result); assert(result ==15566411);
row = 116;
ciphertext_entry =8097162;
#20;
$display("Result = %d", result); assert(result ==8918987);
row = 117;
ciphertext_entry =254588;
#20;
$display("Result = %d", result); assert(result ==11688617);
row = 118;
ciphertext_entry =13211275;
#20;
$display("Result = %d", result); assert(result ==14524575);
row = 119;
ciphertext_entry =5776563;
#20;
$display("Result = %d", result); assert(result ==2303510);
row = 120;
ciphertext_entry =2293504;
#20;
$display("Result = %d", result); assert(result ==14338891);
row = 121;
ciphertext_entry =11126760;
#20;
$display("Result = %d", result); assert(result ==1199734);
row = 122;
ciphertext_entry =2312572;
#20;
$display("Result = %d", result); assert(result ==9089437);
row = 123;
ciphertext_entry =16016002;
#20;
$display("Result = %d", result); assert(result ==10849293);
row = 124;
ciphertext_entry =12841246;
#20;
$display("Result = %d", result); assert(result ==8168630);
row = 125;
ciphertext_entry =7390091;
#20;
$display("Result = %d", result); assert(result ==8814352);
row = 126;
ciphertext_entry =16599182;
#20;
$display("Result = %d", result); assert(result ==6017672);
row = 127;
ciphertext_entry =16668189;
#20;
$display("Result = %d", result); assert(result ==2502774);
row = 128;
ciphertext_entry =1923577;
#20;
$display("Result = %d", result); assert(result ==15497421);
ciphertext_select = 0;
row = 129;
#20;
$display("Result = %d", result); assert(result ==7600909);
row = 130;
#20;
$display("Result = %d", result); assert(result ==4663234);
row = 131;
#20;
$display("Result = %d", result); assert(result ==1642084);
row = 132;
#20;
$display("Result = %d", result); assert(result ==1392776);
row = 133;
#20;
$display("Result = %d", result); assert(result ==1603457);
row = 134;
#20;
$display("Result = %d", result); assert(result ==9124787);
row = 135;
#20;
$display("Result = %d", result); assert(result ==9468087);
row = 136;
#20;
$display("Result = %d", result); assert(result ==14281752);
row = 137;
#20;
$display("Result = %d", result); assert(result ==12975681);
row = 138;
#20;
$display("Result = %d", result); assert(result ==16653978);
row = 139;
#20;
$display("Result = %d", result); assert(result ==13912044);
row = 140;
#20;
$display("Result = %d", result); assert(result ==7550234);
row = 141;
#20;
$display("Result = %d", result); assert(result ==15003264);
row = 142;
#20;
$display("Result = %d", result); assert(result ==16273055);
row = 143;
#20;
$display("Result = %d", result); assert(result ==795857);
row = 144;
#20;
$display("Result = %d", result); assert(result ==6963434);
row = 145;
#20;
$display("Result = %d", result); assert(result ==14451210);
row = 146;
#20;
$display("Result = %d", result); assert(result ==205879);
row = 147;
#20;
$display("Result = %d", result); assert(result ==12773608);
row = 148;
#20;
$display("Result = %d", result); assert(result ==8566451);
row = 149;
#20;
$display("Result = %d", result); assert(result ==12028607);
row = 150;
#20;
$display("Result = %d", result); assert(result ==11485419);
row = 151;
#20;
$display("Result = %d", result); assert(result ==11090266);
row = 152;
#20;
$display("Result = %d", result); assert(result ==3411924);
row = 153;
#20;
$display("Result = %d", result); assert(result ==13012864);
row = 154;
#20;
$display("Result = %d", result); assert(result ==8386698);
row = 155;
#20;
$display("Result = %d", result); assert(result ==3032668);
row = 156;
#20;
$display("Result = %d", result); assert(result ==749900);
row = 157;
#20;
$display("Result = %d", result); assert(result ==4111764);
row = 158;
#20;
$display("Result = %d", result); assert(result ==61346);
row = 159;
#20;
$display("Result = %d", result); assert(result ==9878367);
row = 160;
#20;
$display("Result = %d", result); assert(result ==54492);
row = 161;
#20;
$display("Result = %d", result); assert(result ==7872798);
row = 162;
#20;
$display("Result = %d", result); assert(result ==2583368);
row = 163;
#20;
$display("Result = %d", result); assert(result ==13431394);
row = 164;
#20;
$display("Result = %d", result); assert(result ==1739136);
row = 165;
#20;
$display("Result = %d", result); assert(result ==916642);
row = 166;
#20;
$display("Result = %d", result); assert(result ==6350050);
row = 167;
#20;
$display("Result = %d", result); assert(result ==472141);
row = 168;
#20;
$display("Result = %d", result); assert(result ==2270448);
row = 169;
#20;
$display("Result = %d", result); assert(result ==4426882);
row = 170;
#20;
$display("Result = %d", result); assert(result ==4189681);
row = 171;
#20;
$display("Result = %d", result); assert(result ==7723144);
row = 172;
#20;
$display("Result = %d", result); assert(result ==14831121);
row = 173;
#20;
$display("Result = %d", result); assert(result ==13838354);
row = 174;
#20;
$display("Result = %d", result); assert(result ==8436063);
row = 175;
#20;
$display("Result = %d", result); assert(result ==8370424);
row = 176;
#20;
$display("Result = %d", result); assert(result ==13531415);
row = 177;
#20;
$display("Result = %d", result); assert(result ==6732109);
row = 178;
#20;
$display("Result = %d", result); assert(result ==5784374);
row = 179;
#20;
$display("Result = %d", result); assert(result ==11153093);
row = 180;
#20;
$display("Result = %d", result); assert(result ==14119029);
row = 181;
#20;
$display("Result = %d", result); assert(result ==3020887);
row = 182;
#20;
$display("Result = %d", result); assert(result ==13208682);
row = 183;
#20;
$display("Result = %d", result); assert(result ==1489277);
row = 184;
#20;
$display("Result = %d", result); assert(result ==8320866);
row = 185;
#20;
$display("Result = %d", result); assert(result ==7087915);
row = 186;
#20;
$display("Result = %d", result); assert(result ==13813862);
row = 187;
#20;
$display("Result = %d", result); assert(result ==13470790);
row = 188;
#20;
$display("Result = %d", result); assert(result ==6700896);
row = 189;
#20;
$display("Result = %d", result); assert(result ==2485974);
row = 190;
#20;
$display("Result = %d", result); assert(result ==4967270);
row = 191;
#20;
$display("Result = %d", result); assert(result ==895341);
row = 192;
#20;
$display("Result = %d", result); assert(result ==14263364);
row = 193;
#20;
$display("Result = %d", result); assert(result ==8042125);
row = 194;
#20;
$display("Result = %d", result); assert(result ==16410017);
row = 195;
#20;
$display("Result = %d", result); assert(result ==7065841);
row = 196;
#20;
$display("Result = %d", result); assert(result ==15233309);
row = 197;
#20;
$display("Result = %d", result); assert(result ==8662864);
row = 198;
#20;
$display("Result = %d", result); assert(result ==13987592);
row = 199;
#20;
$display("Result = %d", result); assert(result ==5234494);
row = 200;
#20;
$display("Result = %d", result); assert(result ==3071384);
row = 201;
#20;
$display("Result = %d", result); assert(result ==1839118);
row = 202;
#20;
$display("Result = %d", result); assert(result ==9152437);
row = 203;
#20;
$display("Result = %d", result); assert(result ==10589638);
row = 204;
#20;
$display("Result = %d", result); assert(result ==4819648);
row = 205;
#20;
$display("Result = %d", result); assert(result ==12251436);
row = 206;
#20;
$display("Result = %d", result); assert(result ==9276820);
row = 207;
#20;
$display("Result = %d", result); assert(result ==873390);
row = 208;
#20;
$display("Result = %d", result); assert(result ==12610608);
row = 209;
#20;
$display("Result = %d", result); assert(result ==11941986);
row = 210;
#20;
$display("Result = %d", result); assert(result ==396436);
row = 211;
#20;
$display("Result = %d", result); assert(result ==6489827);
row = 212;
#20;
$display("Result = %d", result); assert(result ==16627110);
row = 213;
#20;
$display("Result = %d", result); assert(result ==10177771);
row = 214;
#20;
$display("Result = %d", result); assert(result ==9604357);
row = 215;
#20;
$display("Result = %d", result); assert(result ==15340521);
row = 216;
#20;
$display("Result = %d", result); assert(result ==4698456);
row = 217;
#20;
$display("Result = %d", result); assert(result ==14109696);
row = 218;
#20;
$display("Result = %d", result); assert(result ==2667151);
row = 219;
#20;
$display("Result = %d", result); assert(result ==10953986);
row = 220;
#20;
$display("Result = %d", result); assert(result ==8808641);
row = 221;
#20;
$display("Result = %d", result); assert(result ==10578529);
row = 222;
#20;
$display("Result = %d", result); assert(result ==14044951);
row = 223;
#20;
$display("Result = %d", result); assert(result ==10023565);
row = 224;
#20;
$display("Result = %d", result); assert(result ==7199366);
row = 225;
#20;
$display("Result = %d", result); assert(result ==16691561);
row = 226;
#20;
$display("Result = %d", result); assert(result ==14793349);
row = 227;
#20;
$display("Result = %d", result); assert(result ==1198060);
row = 228;
#20;
$display("Result = %d", result); assert(result ==2003249);
row = 229;
#20;
$display("Result = %d", result); assert(result ==4720430);
row = 230;
#20;
$display("Result = %d", result); assert(result ==7002262);
row = 231;
#20;
$display("Result = %d", result); assert(result ==7382803);
row = 232;
#20;
$display("Result = %d", result); assert(result ==7736492);
row = 233;
#20;
$display("Result = %d", result); assert(result ==11542101);
row = 234;
#20;
$display("Result = %d", result); assert(result ==12181968);
row = 235;
#20;
$display("Result = %d", result); assert(result ==16372583);
row = 236;
#20;
$display("Result = %d", result); assert(result ==7943846);
row = 237;
#20;
$display("Result = %d", result); assert(result ==12933652);
row = 238;
#20;
$display("Result = %d", result); assert(result ==11547077);
row = 239;
#20;
$display("Result = %d", result); assert(result ==3220871);
row = 240;
#20;
$display("Result = %d", result); assert(result ==4126645);
row = 241;
#20;
$display("Result = %d", result); assert(result ==5704230);
row = 242;
#20;
$display("Result = %d", result); assert(result ==3978646);
row = 243;
#20;
$display("Result = %d", result); assert(result ==6322471);
row = 244;
#20;
$display("Result = %d", result); assert(result ==16320216);
row = 245;
#20;
$display("Result = %d", result); assert(result ==10447999);
row = 246;
#20;
$display("Result = %d", result); assert(result ==4630063);
row = 247;
#20;
$display("Result = %d", result); assert(result ==10254877);
row = 248;
#20;
$display("Result = %d", result); assert(result ==10212492);
row = 249;
#20;
$display("Result = %d", result); assert(result ==15466656);
row = 250;
#20;
$display("Result = %d", result); assert(result ==8660674);
row = 251;
#20;
$display("Result = %d", result); assert(result ==9550370);
row = 252;
#20;
$display("Result = %d", result); assert(result ==12590330);
row = 253;
#20;
$display("Result = %d", result); assert(result ==6125253);
row = 254;
#20;
$display("Result = %d", result); assert(result ==5469706);
row = 255;
#20;
$display("Result = %d", result); assert(result ==10879178);
row = 256;
#20;
$display("Result = %d", result); assert(result ==11523368);
en=0;
rst_n=0;
#100;
rst_n=1;
#100;
en=1;
#20;
ciphertext_select = 0;
row = 0;
ciphertext_entry =3087881;
#20;
row = 1;
ciphertext_entry =4259920;
#20;
row = 2;
ciphertext_entry =11211602;
#20;
row = 3;
ciphertext_entry =14653114;
#20;
row = 4;
ciphertext_entry =15766208;
#20;
row = 5;
ciphertext_entry =14451563;
#20;
row = 6;
ciphertext_entry =5535477;
#20;
row = 7;
ciphertext_entry =15002612;
#20;
row = 8;
ciphertext_entry =14614743;
#20;
row = 9;
ciphertext_entry =9450399;
#20;
row = 10;
ciphertext_entry =4510795;
#20;
row = 11;
ciphertext_entry =912954;
#20;
row = 12;
ciphertext_entry =915869;
#20;
row = 13;
ciphertext_entry =8382521;
#20;
row = 14;
ciphertext_entry =6010876;
#20;
row = 15;
ciphertext_entry =10435820;
#20;
row = 16;
ciphertext_entry =804460;
#20;
row = 17;
ciphertext_entry =528500;
#20;
row = 18;
ciphertext_entry =11380977;
#20;
row = 19;
ciphertext_entry =11523099;
#20;
row = 20;
ciphertext_entry =5709214;
#20;
row = 21;
ciphertext_entry =13496740;
#20;
row = 22;
ciphertext_entry =13778198;
#20;
row = 23;
ciphertext_entry =7628216;
#20;
row = 24;
ciphertext_entry =6136225;
#20;
row = 25;
ciphertext_entry =12997713;
#20;
row = 26;
ciphertext_entry =14582627;
#20;
row = 27;
ciphertext_entry =5130715;
#20;
row = 28;
ciphertext_entry =9809155;
#20;
row = 29;
ciphertext_entry =5811586;
#20;
row = 30;
ciphertext_entry =7073267;
#20;
row = 31;
ciphertext_entry =16162150;
#20;
row = 32;
ciphertext_entry =11144384;
#20;
row = 33;
ciphertext_entry =2617225;
#20;
row = 34;
ciphertext_entry =5398558;
#20;
row = 35;
ciphertext_entry =1229246;
#20;
row = 36;
ciphertext_entry =12484931;
#20;
row = 37;
ciphertext_entry =13764966;
#20;
row = 38;
ciphertext_entry =435501;
#20;
row = 39;
ciphertext_entry =2534371;
#20;
row = 40;
ciphertext_entry =13532297;
#20;
row = 41;
ciphertext_entry =3719937;
#20;
row = 42;
ciphertext_entry =10409516;
#20;
row = 43;
ciphertext_entry =7538322;
#20;
row = 44;
ciphertext_entry =16190767;
#20;
row = 45;
ciphertext_entry =4007760;
#20;
row = 46;
ciphertext_entry =5138873;
#20;
row = 47;
ciphertext_entry =2830729;
#20;
row = 48;
ciphertext_entry =10072731;
#20;
row = 49;
ciphertext_entry =10024961;
#20;
row = 50;
ciphertext_entry =15761992;
#20;
row = 51;
ciphertext_entry =13451076;
#20;
row = 52;
ciphertext_entry =1654891;
#20;
row = 53;
ciphertext_entry =7291603;
#20;
row = 54;
ciphertext_entry =2887190;
#20;
row = 55;
ciphertext_entry =13277339;
#20;
row = 56;
ciphertext_entry =5844243;
#20;
row = 57;
ciphertext_entry =3836430;
#20;
row = 58;
ciphertext_entry =11709160;
#20;
row = 59;
ciphertext_entry =8908558;
#20;
row = 60;
ciphertext_entry =12847668;
#20;
row = 61;
ciphertext_entry =4771138;
#20;
row = 62;
ciphertext_entry =5386695;
#20;
row = 63;
ciphertext_entry =15280239;
#20;
row = 64;
ciphertext_entry =14949715;
#20;
row = 65;
ciphertext_entry =4098460;
#20;
row = 66;
ciphertext_entry =12549220;
#20;
row = 67;
ciphertext_entry =7161052;
#20;
row = 68;
ciphertext_entry =8471115;
#20;
row = 69;
ciphertext_entry =12216823;
#20;
row = 70;
ciphertext_entry =14679941;
#20;
row = 71;
ciphertext_entry =15719535;
#20;
row = 72;
ciphertext_entry =15846075;
#20;
row = 73;
ciphertext_entry =7872181;
#20;
row = 74;
ciphertext_entry =1638804;
#20;
row = 75;
ciphertext_entry =9323396;
#20;
row = 76;
ciphertext_entry =10968666;
#20;
row = 77;
ciphertext_entry =312921;
#20;
row = 78;
ciphertext_entry =398387;
#20;
row = 79;
ciphertext_entry =4198812;
#20;
row = 80;
ciphertext_entry =12799780;
#20;
row = 81;
ciphertext_entry =6756219;
#20;
row = 82;
ciphertext_entry =12946488;
#20;
row = 83;
ciphertext_entry =16602405;
#20;
row = 84;
ciphertext_entry =4905865;
#20;
row = 85;
ciphertext_entry =9115749;
#20;
row = 86;
ciphertext_entry =7408766;
#20;
row = 87;
ciphertext_entry =15442781;
#20;
row = 88;
ciphertext_entry =2759566;
#20;
row = 89;
ciphertext_entry =2000568;
#20;
row = 90;
ciphertext_entry =2176500;
#20;
row = 91;
ciphertext_entry =13014581;
#20;
row = 92;
ciphertext_entry =13188069;
#20;
row = 93;
ciphertext_entry =7115127;
#20;
row = 94;
ciphertext_entry =5028536;
#20;
row = 95;
ciphertext_entry =8583681;
#20;
row = 96;
ciphertext_entry =8431920;
#20;
row = 97;
ciphertext_entry =13458229;
#20;
row = 98;
ciphertext_entry =6550732;
#20;
row = 99;
ciphertext_entry =12158434;
#20;
row = 100;
ciphertext_entry =1324782;
#20;
row = 101;
ciphertext_entry =695627;
#20;
row = 102;
ciphertext_entry =11009740;
#20;
row = 103;
ciphertext_entry =12171714;
#20;
row = 104;
ciphertext_entry =15543099;
#20;
row = 105;
ciphertext_entry =6262300;
#20;
row = 106;
ciphertext_entry =14099345;
#20;
row = 107;
ciphertext_entry =12782151;
#20;
row = 108;
ciphertext_entry =12118365;
#20;
row = 109;
ciphertext_entry =10621042;
#20;
row = 110;
ciphertext_entry =9163321;
#20;
row = 111;
ciphertext_entry =15629871;
#20;
row = 112;
ciphertext_entry =391347;
#20;
row = 113;
ciphertext_entry =3062876;
#20;
row = 114;
ciphertext_entry =33747;
#20;
row = 115;
ciphertext_entry =8089246;
#20;
row = 116;
ciphertext_entry =2309091;
#20;
row = 117;
ciphertext_entry =10339703;
#20;
row = 118;
ciphertext_entry =8542596;
#20;
row = 119;
ciphertext_entry =14549360;
#20;
row = 120;
ciphertext_entry =3626641;
#20;
row = 121;
ciphertext_entry =7666121;
#20;
row = 122;
ciphertext_entry =6712454;
#20;
row = 123;
ciphertext_entry =9713473;
#20;
row = 124;
ciphertext_entry =15205962;
#20;
row = 125;
ciphertext_entry =5174602;
#20;
row = 126;
ciphertext_entry =12059566;
#20;
row = 127;
ciphertext_entry =8594288;
#20;
row = 128;
ciphertext_entry =2197278;
#20;
ciphertext_select = 1;
row = 0;
ciphertext_entry =3087881;
#20;
$display("Result = %d", result); assert(result ==6256294);
row = 1;
ciphertext_entry =4259920;
#20;
$display("Result = %d", result); assert(result ==15131499);
row = 2;
ciphertext_entry =11211602;
#20;
$display("Result = %d", result); assert(result ==16746221);
row = 3;
ciphertext_entry =14653114;
#20;
$display("Result = %d", result); assert(result ==13931842);
row = 4;
ciphertext_entry =15766208;
#20;
$display("Result = %d", result); assert(result ==4407785);
row = 5;
ciphertext_entry =14451563;
#20;
$display("Result = %d", result); assert(result ==7186238);
row = 6;
ciphertext_entry =5535477;
#20;
$display("Result = %d", result); assert(result ==3688615);
row = 7;
ciphertext_entry =15002612;
#20;
$display("Result = %d", result); assert(result ==10666035);
row = 8;
ciphertext_entry =14614743;
#20;
$display("Result = %d", result); assert(result ==685167);
row = 9;
ciphertext_entry =9450399;
#20;
$display("Result = %d", result); assert(result ==1161987);
row = 10;
ciphertext_entry =4510795;
#20;
$display("Result = %d", result); assert(result ==7440584);
row = 11;
ciphertext_entry =912954;
#20;
$display("Result = %d", result); assert(result ==15971410);
row = 12;
ciphertext_entry =915869;
#20;
$display("Result = %d", result); assert(result ==6514308);
row = 13;
ciphertext_entry =8382521;
#20;
$display("Result = %d", result); assert(result ==7508077);
row = 14;
ciphertext_entry =6010876;
#20;
$display("Result = %d", result); assert(result ==11621683);
row = 15;
ciphertext_entry =10435820;
#20;
$display("Result = %d", result); assert(result ==12434905);
row = 16;
ciphertext_entry =804460;
#20;
$display("Result = %d", result); assert(result ==8355498);
row = 17;
ciphertext_entry =528500;
#20;
$display("Result = %d", result); assert(result ==15218846);
row = 18;
ciphertext_entry =11380977;
#20;
$display("Result = %d", result); assert(result ==14583794);
row = 19;
ciphertext_entry =11523099;
#20;
$display("Result = %d", result); assert(result ==4555924);
row = 20;
ciphertext_entry =5709214;
#20;
$display("Result = %d", result); assert(result ==794642);
row = 21;
ciphertext_entry =13496740;
#20;
$display("Result = %d", result); assert(result ==10187240);
row = 22;
ciphertext_entry =13778198;
#20;
$display("Result = %d", result); assert(result ==10923964);
row = 23;
ciphertext_entry =7628216;
#20;
$display("Result = %d", result); assert(result ==8389382);
row = 24;
ciphertext_entry =6136225;
#20;
$display("Result = %d", result); assert(result ==4210938);
row = 25;
ciphertext_entry =12997713;
#20;
$display("Result = %d", result); assert(result ==119949);
row = 26;
ciphertext_entry =14582627;
#20;
$display("Result = %d", result); assert(result ==7700149);
row = 27;
ciphertext_entry =5130715;
#20;
$display("Result = %d", result); assert(result ==7864993);
row = 28;
ciphertext_entry =9809155;
#20;
$display("Result = %d", result); assert(result ==13805601);
row = 29;
ciphertext_entry =5811586;
#20;
$display("Result = %d", result); assert(result ==2821079);
row = 30;
ciphertext_entry =7073267;
#20;
$display("Result = %d", result); assert(result ==16096454);
row = 31;
ciphertext_entry =16162150;
#20;
$display("Result = %d", result); assert(result ==5343952);
row = 32;
ciphertext_entry =11144384;
#20;
$display("Result = %d", result); assert(result ==16142251);
row = 33;
ciphertext_entry =2617225;
#20;
$display("Result = %d", result); assert(result ==10461883);
row = 34;
ciphertext_entry =5398558;
#20;
$display("Result = %d", result); assert(result ==10774025);
row = 35;
ciphertext_entry =1229246;
#20;
$display("Result = %d", result); assert(result ==5892439);
row = 36;
ciphertext_entry =12484931;
#20;
$display("Result = %d", result); assert(result ==14414970);
row = 37;
ciphertext_entry =13764966;
#20;
$display("Result = %d", result); assert(result ==8741432);
row = 38;
ciphertext_entry =435501;
#20;
$display("Result = %d", result); assert(result ==13611712);
row = 39;
ciphertext_entry =2534371;
#20;
$display("Result = %d", result); assert(result ==10382345);
row = 40;
ciphertext_entry =13532297;
#20;
$display("Result = %d", result); assert(result ==5133261);
row = 41;
ciphertext_entry =3719937;
#20;
$display("Result = %d", result); assert(result ==10987807);
row = 42;
ciphertext_entry =10409516;
#20;
$display("Result = %d", result); assert(result ==13395716);
row = 43;
ciphertext_entry =7538322;
#20;
$display("Result = %d", result); assert(result ==14489586);
row = 44;
ciphertext_entry =16190767;
#20;
$display("Result = %d", result); assert(result ==516668);
row = 45;
ciphertext_entry =4007760;
#20;
$display("Result = %d", result); assert(result ==8146030);
row = 46;
ciphertext_entry =5138873;
#20;
$display("Result = %d", result); assert(result ==1767921);
row = 47;
ciphertext_entry =2830729;
#20;
$display("Result = %d", result); assert(result ==8068794);
row = 48;
ciphertext_entry =10072731;
#20;
$display("Result = %d", result); assert(result ==5145410);
row = 49;
ciphertext_entry =10024961;
#20;
$display("Result = %d", result); assert(result ==6124160);
row = 50;
ciphertext_entry =15761992;
#20;
$display("Result = %d", result); assert(result ==2539287);
row = 51;
ciphertext_entry =13451076;
#20;
$display("Result = %d", result); assert(result ==3405589);
row = 52;
ciphertext_entry =1654891;
#20;
$display("Result = %d", result); assert(result ==10212585);
row = 53;
ciphertext_entry =7291603;
#20;
$display("Result = %d", result); assert(result ==15757449);
row = 54;
ciphertext_entry =2887190;
#20;
$display("Result = %d", result); assert(result ==7322616);
row = 55;
ciphertext_entry =13277339;
#20;
$display("Result = %d", result); assert(result ==9539706);
row = 56;
ciphertext_entry =5844243;
#20;
$display("Result = %d", result); assert(result ==1237883);
row = 57;
ciphertext_entry =3836430;
#20;
$display("Result = %d", result); assert(result ==2459214);
row = 58;
ciphertext_entry =11709160;
#20;
$display("Result = %d", result); assert(result ==2472279);
row = 59;
ciphertext_entry =8908558;
#20;
$display("Result = %d", result); assert(result ==15269789);
row = 60;
ciphertext_entry =12847668;
#20;
$display("Result = %d", result); assert(result ==698077);
row = 61;
ciphertext_entry =4771138;
#20;
$display("Result = %d", result); assert(result ==16414170);
row = 62;
ciphertext_entry =5386695;
#20;
$display("Result = %d", result); assert(result ==6288182);
row = 63;
ciphertext_entry =15280239;
#20;
$display("Result = %d", result); assert(result ==11101629);
row = 64;
ciphertext_entry =14949715;
#20;
$display("Result = %d", result); assert(result ==16341874);
row = 65;
ciphertext_entry =4098460;
#20;
$display("Result = %d", result); assert(result ==14887629);
row = 66;
ciphertext_entry =12549220;
#20;
$display("Result = %d", result); assert(result ==14891512);
row = 67;
ciphertext_entry =7161052;
#20;
$display("Result = %d", result); assert(result ==16520800);
row = 68;
ciphertext_entry =8471115;
#20;
$display("Result = %d", result); assert(result ==4746515);
row = 69;
ciphertext_entry =12216823;
#20;
$display("Result = %d", result); assert(result ==9273872);
row = 70;
ciphertext_entry =14679941;
#20;
$display("Result = %d", result); assert(result ==14091068);
row = 71;
ciphertext_entry =15719535;
#20;
$display("Result = %d", result); assert(result ==16229309);
row = 72;
ciphertext_entry =15846075;
#20;
$display("Result = %d", result); assert(result ==13850498);
row = 73;
ciphertext_entry =7872181;
#20;
$display("Result = %d", result); assert(result ==10285814);
row = 74;
ciphertext_entry =1638804;
#20;
$display("Result = %d", result); assert(result ==791127);
row = 75;
ciphertext_entry =9323396;
#20;
$display("Result = %d", result); assert(result ==5711425);
row = 76;
ciphertext_entry =10968666;
#20;
$display("Result = %d", result); assert(result ==1111543);
row = 77;
ciphertext_entry =312921;
#20;
$display("Result = %d", result); assert(result ==9722806);
row = 78;
ciphertext_entry =398387;
#20;
$display("Result = %d", result); assert(result ==2542199);
row = 79;
ciphertext_entry =4198812;
#20;
$display("Result = %d", result); assert(result ==272633);
row = 80;
ciphertext_entry =12799780;
#20;
$display("Result = %d", result); assert(result ==14875797);
row = 81;
ciphertext_entry =6756219;
#20;
$display("Result = %d", result); assert(result ==16039321);
row = 82;
ciphertext_entry =12946488;
#20;
$display("Result = %d", result); assert(result ==4453264);
row = 83;
ciphertext_entry =16602405;
#20;
$display("Result = %d", result); assert(result ==14237665);
row = 84;
ciphertext_entry =4905865;
#20;
$display("Result = %d", result); assert(result ==3379915);
row = 85;
ciphertext_entry =9115749;
#20;
$display("Result = %d", result); assert(result ==775013);
row = 86;
ciphertext_entry =7408766;
#20;
$display("Result = %d", result); assert(result ==16205038);
row = 87;
ciphertext_entry =15442781;
#20;
$display("Result = %d", result); assert(result ==4386753);
row = 88;
ciphertext_entry =2759566;
#20;
$display("Result = %d", result); assert(result ==1549595);
row = 89;
ciphertext_entry =2000568;
#20;
$display("Result = %d", result); assert(result ==3026444);
row = 90;
ciphertext_entry =2176500;
#20;
$display("Result = %d", result); assert(result ==8442575);
row = 91;
ciphertext_entry =13014581;
#20;
$display("Result = %d", result); assert(result ==9366125);
row = 92;
ciphertext_entry =13188069;
#20;
$display("Result = %d", result); assert(result ==16294380);
row = 93;
ciphertext_entry =7115127;
#20;
$display("Result = %d", result); assert(result ==12431523);
row = 94;
ciphertext_entry =5028536;
#20;
$display("Result = %d", result); assert(result ==16358453);
row = 95;
ciphertext_entry =8583681;
#20;
$display("Result = %d", result); assert(result ==11200461);
row = 96;
ciphertext_entry =8431920;
#20;
$display("Result = %d", result); assert(result ==2346168);
row = 97;
ciphertext_entry =13458229;
#20;
$display("Result = %d", result); assert(result ==4329614);
row = 98;
ciphertext_entry =6550732;
#20;
$display("Result = %d", result); assert(result ==10358430);
row = 99;
ciphertext_entry =12158434;
#20;
$display("Result = %d", result); assert(result ==4096634);
row = 100;
ciphertext_entry =1324782;
#20;
$display("Result = %d", result); assert(result ==16390328);
row = 101;
ciphertext_entry =695627;
#20;
$display("Result = %d", result); assert(result ==8966616);
row = 102;
ciphertext_entry =11009740;
#20;
$display("Result = %d", result); assert(result ==6881415);
row = 103;
ciphertext_entry =12171714;
#20;
$display("Result = %d", result); assert(result ==1376132);
row = 104;
ciphertext_entry =15543099;
#20;
$display("Result = %d", result); assert(result ==11882793);
row = 105;
ciphertext_entry =6262300;
#20;
$display("Result = %d", result); assert(result ==15542983);
row = 106;
ciphertext_entry =14099345;
#20;
$display("Result = %d", result); assert(result ==13240093);
row = 107;
ciphertext_entry =12782151;
#20;
$display("Result = %d", result); assert(result ==1555293);
row = 108;
ciphertext_entry =12118365;
#20;
$display("Result = %d", result); assert(result ==10501641);
row = 109;
ciphertext_entry =10621042;
#20;
$display("Result = %d", result); assert(result ==11554665);
row = 110;
ciphertext_entry =9163321;
#20;
$display("Result = %d", result); assert(result ==9488632);
row = 111;
ciphertext_entry =15629871;
#20;
$display("Result = %d", result); assert(result ==14171716);
row = 112;
ciphertext_entry =391347;
#20;
$display("Result = %d", result); assert(result ==1331473);
row = 113;
ciphertext_entry =3062876;
#20;
$display("Result = %d", result); assert(result ==888694);
row = 114;
ciphertext_entry =33747;
#20;
$display("Result = %d", result); assert(result ==7131516);
row = 115;
ciphertext_entry =8089246;
#20;
$display("Result = %d", result); assert(result ==6960453);
row = 116;
ciphertext_entry =2309091;
#20;
$display("Result = %d", result); assert(result ==9703713);
row = 117;
ciphertext_entry =10339703;
#20;
$display("Result = %d", result); assert(result ==8053682);
row = 118;
ciphertext_entry =8542596;
#20;
$display("Result = %d", result); assert(result ==13320316);
row = 119;
ciphertext_entry =14549360;
#20;
$display("Result = %d", result); assert(result ==15994752);
row = 120;
ciphertext_entry =3626641;
#20;
$display("Result = %d", result); assert(result ==4376390);
row = 121;
ciphertext_entry =7666121;
#20;
$display("Result = %d", result); assert(result ==11869365);
row = 122;
ciphertext_entry =6712454;
#20;
$display("Result = %d", result); assert(result ==10917546);
row = 123;
ciphertext_entry =9713473;
#20;
$display("Result = %d", result); assert(result ==16195737);
row = 124;
ciphertext_entry =15205962;
#20;
$display("Result = %d", result); assert(result ==7141126);
row = 125;
ciphertext_entry =5174602;
#20;
$display("Result = %d", result); assert(result ==6548602);
row = 126;
ciphertext_entry =12059566;
#20;
$display("Result = %d", result); assert(result ==12422764);
row = 127;
ciphertext_entry =8594288;
#20;
$display("Result = %d", result); assert(result ==13311150);
row = 128;
ciphertext_entry =2197278;
#20;
$display("Result = %d", result); assert(result ==8252750);
ciphertext_select = 0;
row = 129;
#20;
$display("Result = %d", result); assert(result ==2463568);
row = 130;
#20;
$display("Result = %d", result); assert(result ==15720963);
row = 131;
#20;
$display("Result = %d", result); assert(result ==2171679);
row = 132;
#20;
$display("Result = %d", result); assert(result ==12901611);
row = 133;
#20;
$display("Result = %d", result); assert(result ==2304686);
row = 134;
#20;
$display("Result = %d", result); assert(result ==11589821);
row = 135;
#20;
$display("Result = %d", result); assert(result ==14809958);
row = 136;
#20;
$display("Result = %d", result); assert(result ==6003673);
row = 137;
#20;
$display("Result = %d", result); assert(result ==3900575);
row = 138;
#20;
$display("Result = %d", result); assert(result ==7596275);
row = 139;
#20;
$display("Result = %d", result); assert(result ==7235363);
row = 140;
#20;
$display("Result = %d", result); assert(result ==13549652);
row = 141;
#20;
$display("Result = %d", result); assert(result ==15573153);
row = 142;
#20;
$display("Result = %d", result); assert(result ==408824);
row = 143;
#20;
$display("Result = %d", result); assert(result ==7276653);
row = 144;
#20;
$display("Result = %d", result); assert(result ==11367527);
row = 145;
#20;
$display("Result = %d", result); assert(result ==12798301);
row = 146;
#20;
$display("Result = %d", result); assert(result ==16599335);
row = 147;
#20;
$display("Result = %d", result); assert(result ==9635923);
row = 148;
#20;
$display("Result = %d", result); assert(result ==853925);
row = 149;
#20;
$display("Result = %d", result); assert(result ==4160099);
row = 150;
#20;
$display("Result = %d", result); assert(result ==16447799);
row = 151;
#20;
$display("Result = %d", result); assert(result ==2911215);
row = 152;
#20;
$display("Result = %d", result); assert(result ==13502832);
row = 153;
#20;
$display("Result = %d", result); assert(result ==10391880);
row = 154;
#20;
$display("Result = %d", result); assert(result ==10961699);
row = 155;
#20;
$display("Result = %d", result); assert(result ==3629361);
row = 156;
#20;
$display("Result = %d", result); assert(result ==6889534);
row = 157;
#20;
$display("Result = %d", result); assert(result ==4340743);
row = 158;
#20;
$display("Result = %d", result); assert(result ==15723555);
row = 159;
#20;
$display("Result = %d", result); assert(result ==3362354);
row = 160;
#20;
$display("Result = %d", result); assert(result ==3007670);
row = 161;
#20;
$display("Result = %d", result); assert(result ==10277154);
row = 162;
#20;
$display("Result = %d", result); assert(result ==14487843);
row = 163;
#20;
$display("Result = %d", result); assert(result ==10600755);
row = 164;
#20;
$display("Result = %d", result); assert(result ==11821690);
row = 165;
#20;
$display("Result = %d", result); assert(result ==3647719);
row = 166;
#20;
$display("Result = %d", result); assert(result ==4989155);
row = 167;
#20;
$display("Result = %d", result); assert(result ==3667771);
row = 168;
#20;
$display("Result = %d", result); assert(result ==8345033);
row = 169;
#20;
$display("Result = %d", result); assert(result ==5693591);
row = 170;
#20;
$display("Result = %d", result); assert(result ==1516956);
row = 171;
#20;
$display("Result = %d", result); assert(result ==1958366);
row = 172;
#20;
$display("Result = %d", result); assert(result ==443001);
row = 173;
#20;
$display("Result = %d", result); assert(result ==9945917);
row = 174;
#20;
$display("Result = %d", result); assert(result ==10387567);
row = 175;
#20;
$display("Result = %d", result); assert(result ==8515980);
row = 176;
#20;
$display("Result = %d", result); assert(result ==12580124);
row = 177;
#20;
$display("Result = %d", result); assert(result ==9415605);
row = 178;
#20;
$display("Result = %d", result); assert(result ==12997305);
row = 179;
#20;
$display("Result = %d", result); assert(result ==5544733);
row = 180;
#20;
$display("Result = %d", result); assert(result ==6670928);
row = 181;
#20;
$display("Result = %d", result); assert(result ==1627438);
row = 182;
#20;
$display("Result = %d", result); assert(result ==290518);
row = 183;
#20;
$display("Result = %d", result); assert(result ==7726627);
row = 184;
#20;
$display("Result = %d", result); assert(result ==4988749);
row = 185;
#20;
$display("Result = %d", result); assert(result ==14196892);
row = 186;
#20;
$display("Result = %d", result); assert(result ==6487416);
row = 187;
#20;
$display("Result = %d", result); assert(result ==11353620);
row = 188;
#20;
$display("Result = %d", result); assert(result ==4946113);
row = 189;
#20;
$display("Result = %d", result); assert(result ==8188522);
row = 190;
#20;
$display("Result = %d", result); assert(result ==5638849);
row = 191;
#20;
$display("Result = %d", result); assert(result ==7134211);
row = 192;
#20;
$display("Result = %d", result); assert(result ==7001974);
row = 193;
#20;
$display("Result = %d", result); assert(result ==5485599);
row = 194;
#20;
$display("Result = %d", result); assert(result ==3480242);
row = 195;
#20;
$display("Result = %d", result); assert(result ==14341840);
row = 196;
#20;
$display("Result = %d", result); assert(result ==3899209);
row = 197;
#20;
$display("Result = %d", result); assert(result ==9820551);
row = 198;
#20;
$display("Result = %d", result); assert(result ==15261271);
row = 199;
#20;
$display("Result = %d", result); assert(result ==5767675);
row = 200;
#20;
$display("Result = %d", result); assert(result ==16653462);
row = 201;
#20;
$display("Result = %d", result); assert(result ==999307);
row = 202;
#20;
$display("Result = %d", result); assert(result ==15156191);
row = 203;
#20;
$display("Result = %d", result); assert(result ==12764430);
row = 204;
#20;
$display("Result = %d", result); assert(result ==13050816);
row = 205;
#20;
$display("Result = %d", result); assert(result ==6038872);
row = 206;
#20;
$display("Result = %d", result); assert(result ==12193247);
row = 207;
#20;
$display("Result = %d", result); assert(result ==14764451);
row = 208;
#20;
$display("Result = %d", result); assert(result ==6804321);
row = 209;
#20;
$display("Result = %d", result); assert(result ==2923664);
row = 210;
#20;
$display("Result = %d", result); assert(result ==9769429);
row = 211;
#20;
$display("Result = %d", result); assert(result ==13710048);
row = 212;
#20;
$display("Result = %d", result); assert(result ==14135390);
row = 213;
#20;
$display("Result = %d", result); assert(result ==11031932);
row = 214;
#20;
$display("Result = %d", result); assert(result ==10265764);
row = 215;
#20;
$display("Result = %d", result); assert(result ==9396780);
row = 216;
#20;
$display("Result = %d", result); assert(result ==7126977);
row = 217;
#20;
$display("Result = %d", result); assert(result ==1184870);
row = 218;
#20;
$display("Result = %d", result); assert(result ==6069395);
row = 219;
#20;
$display("Result = %d", result); assert(result ==11095595);
row = 220;
#20;
$display("Result = %d", result); assert(result ==12926424);
row = 221;
#20;
$display("Result = %d", result); assert(result ==11201451);
row = 222;
#20;
$display("Result = %d", result); assert(result ==12562742);
row = 223;
#20;
$display("Result = %d", result); assert(result ==16606147);
row = 224;
#20;
$display("Result = %d", result); assert(result ==5881194);
row = 225;
#20;
$display("Result = %d", result); assert(result ==5059241);
row = 226;
#20;
$display("Result = %d", result); assert(result ==11289064);
row = 227;
#20;
$display("Result = %d", result); assert(result ==5120958);
row = 228;
#20;
$display("Result = %d", result); assert(result ==13717045);
row = 229;
#20;
$display("Result = %d", result); assert(result ==8942091);
row = 230;
#20;
$display("Result = %d", result); assert(result ==1579911);
row = 231;
#20;
$display("Result = %d", result); assert(result ==3772551);
row = 232;
#20;
$display("Result = %d", result); assert(result ==6004922);
row = 233;
#20;
$display("Result = %d", result); assert(result ==5505784);
row = 234;
#20;
$display("Result = %d", result); assert(result ==5379803);
row = 235;
#20;
$display("Result = %d", result); assert(result ==9450707);
row = 236;
#20;
$display("Result = %d", result); assert(result ==2743001);
row = 237;
#20;
$display("Result = %d", result); assert(result ==1226000);
row = 238;
#20;
$display("Result = %d", result); assert(result ==14593061);
row = 239;
#20;
$display("Result = %d", result); assert(result ==2497783);
row = 240;
#20;
$display("Result = %d", result); assert(result ==8535391);
row = 241;
#20;
$display("Result = %d", result); assert(result ==9998764);
row = 242;
#20;
$display("Result = %d", result); assert(result ==11279748);
row = 243;
#20;
$display("Result = %d", result); assert(result ==14989547);
row = 244;
#20;
$display("Result = %d", result); assert(result ==15373422);
row = 245;
#20;
$display("Result = %d", result); assert(result ==14262089);
row = 246;
#20;
$display("Result = %d", result); assert(result ==9091975);
row = 247;
#20;
$display("Result = %d", result); assert(result ==12879122);
row = 248;
#20;
$display("Result = %d", result); assert(result ==1134078);
row = 249;
#20;
$display("Result = %d", result); assert(result ==13934080);
row = 250;
#20;
$display("Result = %d", result); assert(result ==9129169);
row = 251;
#20;
$display("Result = %d", result); assert(result ==3279708);
row = 252;
#20;
$display("Result = %d", result); assert(result ==8394216);
row = 253;
#20;
$display("Result = %d", result); assert(result ==9440496);
row = 254;
#20;
$display("Result = %d", result); assert(result ==16310268);
row = 255;
#20;
$display("Result = %d", result); assert(result ==6998538);
row = 256;
#20;
$display("Result = %d", result); assert(result ==13728448);

$finish;
end
endmodule
            
