`define PLAINTEXT_MODULUS 32
`define PLAINTEXT_WIDTH 5
`define DIMENSION 128
`define CIPHERTEXT_MODULUS 16777216
`define CIPHERTEXT_WIDTH 24
`define BIG_N 6425

module decrypt_tb;

    reg clk;
    reg rst_n;
    reg [`CIPHERTEXT_WIDTH-1:0] secret_key [`DIMENSION:0];
    reg signed [`CIPHERTEXT_WIDTH-1:0] cipher_text [`DIMENSION:0];
    reg [`CIPHERTEXT_WIDTH-1:0] skentry;
    reg signed [`CIPHERTEXT_WIDTH-1:0] ctentry;
    reg [`DIMENSION:0] row;
    wire [`PLAINTEXT_WIDTH-1:0] result;
    reg [`PLAINTEXT_WIDTH-1:0] expected;

    always #10 clk = ~clk;

    decrypt #(
        .PLAINTEXT_MODULUS(`PLAINTEXT_MODULUS),
        .PLAINTEXT_WIDTH(`PLAINTEXT_WIDTH),
        .CIPHERTEXT_MODULUS(`CIPHERTEXT_MODULUS),
        .CIPHERTEXT_WIDTH(`CIPHERTEXT_WIDTH),
        .DIMENSION(`DIMENSION),
        .BIG_N(`BIG_N)
    ) decrypt_inst (
        .clk(clk),
        .rst_n(rst_n),
        .secretkey_entry(skentry),
        .ciphertext_entry(ctentry),
        .row(row),
        .result(result)
    );

    initial begin

secret_key[0] = `CIPHERTEXT_WIDTH'd1;
secret_key[1] = `CIPHERTEXT_WIDTH'd2914804;
secret_key[2] = `CIPHERTEXT_WIDTH'd7111320;
secret_key[3] = `CIPHERTEXT_WIDTH'd9764306;
secret_key[4] = `CIPHERTEXT_WIDTH'd16270169;
secret_key[5] = `CIPHERTEXT_WIDTH'd2477246;
secret_key[6] = `CIPHERTEXT_WIDTH'd2470477;
secret_key[7] = `CIPHERTEXT_WIDTH'd7233846;
secret_key[8] = `CIPHERTEXT_WIDTH'd7622992;
secret_key[9] = `CIPHERTEXT_WIDTH'd10474204;
secret_key[10] = `CIPHERTEXT_WIDTH'd9180602;
secret_key[11] = `CIPHERTEXT_WIDTH'd13868973;
secret_key[12] = `CIPHERTEXT_WIDTH'd6779138;
secret_key[13] = `CIPHERTEXT_WIDTH'd9718670;
secret_key[14] = `CIPHERTEXT_WIDTH'd8876301;
secret_key[15] = `CIPHERTEXT_WIDTH'd3219549;
secret_key[16] = `CIPHERTEXT_WIDTH'd6544466;
secret_key[17] = `CIPHERTEXT_WIDTH'd4772816;
secret_key[18] = `CIPHERTEXT_WIDTH'd15806570;
secret_key[19] = `CIPHERTEXT_WIDTH'd10947635;
secret_key[20] = `CIPHERTEXT_WIDTH'd4167960;
secret_key[21] = `CIPHERTEXT_WIDTH'd8438746;
secret_key[22] = `CIPHERTEXT_WIDTH'd12676654;
secret_key[23] = `CIPHERTEXT_WIDTH'd1272369;
secret_key[24] = `CIPHERTEXT_WIDTH'd7862804;
secret_key[25] = `CIPHERTEXT_WIDTH'd9571549;
secret_key[26] = `CIPHERTEXT_WIDTH'd4201878;
secret_key[27] = `CIPHERTEXT_WIDTH'd6873582;
secret_key[28] = `CIPHERTEXT_WIDTH'd7860835;
secret_key[29] = `CIPHERTEXT_WIDTH'd6991297;
secret_key[30] = `CIPHERTEXT_WIDTH'd1151011;
secret_key[31] = `CIPHERTEXT_WIDTH'd5342226;
secret_key[32] = `CIPHERTEXT_WIDTH'd15118860;
secret_key[33] = `CIPHERTEXT_WIDTH'd13466507;
secret_key[34] = `CIPHERTEXT_WIDTH'd14228721;
secret_key[35] = `CIPHERTEXT_WIDTH'd4921273;
secret_key[36] = `CIPHERTEXT_WIDTH'd425177;
secret_key[37] = `CIPHERTEXT_WIDTH'd10620987;
secret_key[38] = `CIPHERTEXT_WIDTH'd5285133;
secret_key[39] = `CIPHERTEXT_WIDTH'd13368943;
secret_key[40] = `CIPHERTEXT_WIDTH'd8664412;
secret_key[41] = `CIPHERTEXT_WIDTH'd4607069;
secret_key[42] = `CIPHERTEXT_WIDTH'd3702434;
secret_key[43] = `CIPHERTEXT_WIDTH'd13683025;
secret_key[44] = `CIPHERTEXT_WIDTH'd7130923;
secret_key[45] = `CIPHERTEXT_WIDTH'd12081749;
secret_key[46] = `CIPHERTEXT_WIDTH'd12079787;
secret_key[47] = `CIPHERTEXT_WIDTH'd4960906;
secret_key[48] = `CIPHERTEXT_WIDTH'd16390017;
secret_key[49] = `CIPHERTEXT_WIDTH'd3115058;
secret_key[50] = `CIPHERTEXT_WIDTH'd3402892;
secret_key[51] = `CIPHERTEXT_WIDTH'd14322125;
secret_key[52] = `CIPHERTEXT_WIDTH'd11805533;
secret_key[53] = `CIPHERTEXT_WIDTH'd7656929;
secret_key[54] = `CIPHERTEXT_WIDTH'd7389158;
secret_key[55] = `CIPHERTEXT_WIDTH'd15104642;
secret_key[56] = `CIPHERTEXT_WIDTH'd16580716;
secret_key[57] = `CIPHERTEXT_WIDTH'd8932987;
secret_key[58] = `CIPHERTEXT_WIDTH'd1735861;
secret_key[59] = `CIPHERTEXT_WIDTH'd5858510;
secret_key[60] = `CIPHERTEXT_WIDTH'd11357771;
secret_key[61] = `CIPHERTEXT_WIDTH'd15726598;
secret_key[62] = `CIPHERTEXT_WIDTH'd13642483;
secret_key[63] = `CIPHERTEXT_WIDTH'd3305697;
secret_key[64] = `CIPHERTEXT_WIDTH'd9758396;
secret_key[65] = `CIPHERTEXT_WIDTH'd5220598;
secret_key[66] = `CIPHERTEXT_WIDTH'd1342696;
secret_key[67] = `CIPHERTEXT_WIDTH'd12243828;
secret_key[68] = `CIPHERTEXT_WIDTH'd12508842;
secret_key[69] = `CIPHERTEXT_WIDTH'd2088854;
secret_key[70] = `CIPHERTEXT_WIDTH'd16123863;
secret_key[71] = `CIPHERTEXT_WIDTH'd14850853;
secret_key[72] = `CIPHERTEXT_WIDTH'd14138285;
secret_key[73] = `CIPHERTEXT_WIDTH'd4711052;
secret_key[74] = `CIPHERTEXT_WIDTH'd15553693;
secret_key[75] = `CIPHERTEXT_WIDTH'd4451789;
secret_key[76] = `CIPHERTEXT_WIDTH'd530002;
secret_key[77] = `CIPHERTEXT_WIDTH'd2564492;
secret_key[78] = `CIPHERTEXT_WIDTH'd10197680;
secret_key[79] = `CIPHERTEXT_WIDTH'd9612489;
secret_key[80] = `CIPHERTEXT_WIDTH'd9957003;
secret_key[81] = `CIPHERTEXT_WIDTH'd13716290;
secret_key[82] = `CIPHERTEXT_WIDTH'd16733561;
secret_key[83] = `CIPHERTEXT_WIDTH'd10775786;
secret_key[84] = `CIPHERTEXT_WIDTH'd2264105;
secret_key[85] = `CIPHERTEXT_WIDTH'd15716264;
secret_key[86] = `CIPHERTEXT_WIDTH'd11583145;
secret_key[87] = `CIPHERTEXT_WIDTH'd4710457;
secret_key[88] = `CIPHERTEXT_WIDTH'd13889942;
secret_key[89] = `CIPHERTEXT_WIDTH'd621457;
secret_key[90] = `CIPHERTEXT_WIDTH'd12416167;
secret_key[91] = `CIPHERTEXT_WIDTH'd10282098;
secret_key[92] = `CIPHERTEXT_WIDTH'd11969588;
secret_key[93] = `CIPHERTEXT_WIDTH'd16242934;
secret_key[94] = `CIPHERTEXT_WIDTH'd5894750;
secret_key[95] = `CIPHERTEXT_WIDTH'd2757712;
secret_key[96] = `CIPHERTEXT_WIDTH'd11787413;
secret_key[97] = `CIPHERTEXT_WIDTH'd13790505;
secret_key[98] = `CIPHERTEXT_WIDTH'd7024878;
secret_key[99] = `CIPHERTEXT_WIDTH'd9628723;
secret_key[100] = `CIPHERTEXT_WIDTH'd12637654;
secret_key[101] = `CIPHERTEXT_WIDTH'd3168378;
secret_key[102] = `CIPHERTEXT_WIDTH'd12781480;
secret_key[103] = `CIPHERTEXT_WIDTH'd15111488;
secret_key[104] = `CIPHERTEXT_WIDTH'd16585117;
secret_key[105] = `CIPHERTEXT_WIDTH'd6075920;
secret_key[106] = `CIPHERTEXT_WIDTH'd14591473;
secret_key[107] = `CIPHERTEXT_WIDTH'd6287864;
secret_key[108] = `CIPHERTEXT_WIDTH'd10320466;
secret_key[109] = `CIPHERTEXT_WIDTH'd10833124;
secret_key[110] = `CIPHERTEXT_WIDTH'd11989945;
secret_key[111] = `CIPHERTEXT_WIDTH'd4255908;
secret_key[112] = `CIPHERTEXT_WIDTH'd9438919;
secret_key[113] = `CIPHERTEXT_WIDTH'd12149259;
secret_key[114] = `CIPHERTEXT_WIDTH'd9735961;
secret_key[115] = `CIPHERTEXT_WIDTH'd1922428;
secret_key[116] = `CIPHERTEXT_WIDTH'd16264759;
secret_key[117] = `CIPHERTEXT_WIDTH'd5909865;
secret_key[118] = `CIPHERTEXT_WIDTH'd11089605;
secret_key[119] = `CIPHERTEXT_WIDTH'd3571527;
secret_key[120] = `CIPHERTEXT_WIDTH'd6333540;
secret_key[121] = `CIPHERTEXT_WIDTH'd9139546;
secret_key[122] = `CIPHERTEXT_WIDTH'd3439654;
secret_key[123] = `CIPHERTEXT_WIDTH'd16320988;
secret_key[124] = `CIPHERTEXT_WIDTH'd3260666;
secret_key[125] = `CIPHERTEXT_WIDTH'd6940522;
secret_key[126] = `CIPHERTEXT_WIDTH'd14190365;
secret_key[127] = `CIPHERTEXT_WIDTH'd16189298;
expected = 0;
cipher_text[0] = `CIPHERTEXT_WIDTH'd11878251;
cipher_text[1] = `CIPHERTEXT_WIDTH'd391936;
cipher_text[2] = `CIPHERTEXT_WIDTH'd8239380;
cipher_text[3] = `CIPHERTEXT_WIDTH'd5863366;
cipher_text[4] = `CIPHERTEXT_WIDTH'd13626513;
cipher_text[5] = `CIPHERTEXT_WIDTH'd4860891;
cipher_text[6] = `CIPHERTEXT_WIDTH'd5351503;
cipher_text[7] = `CIPHERTEXT_WIDTH'd16643855;
cipher_text[8] = `CIPHERTEXT_WIDTH'd1104138;
cipher_text[9] = `CIPHERTEXT_WIDTH'd3493932;
cipher_text[10] = `CIPHERTEXT_WIDTH'd2674594;
cipher_text[11] = `CIPHERTEXT_WIDTH'd7985843;
cipher_text[12] = `CIPHERTEXT_WIDTH'd10531735;
cipher_text[13] = `CIPHERTEXT_WIDTH'd5573010;
cipher_text[14] = `CIPHERTEXT_WIDTH'd4912605;
cipher_text[15] = `CIPHERTEXT_WIDTH'd8262899;
cipher_text[16] = `CIPHERTEXT_WIDTH'd16646916;
cipher_text[17] = `CIPHERTEXT_WIDTH'd14381706;
cipher_text[18] = `CIPHERTEXT_WIDTH'd12297390;
cipher_text[19] = `CIPHERTEXT_WIDTH'd13413363;
cipher_text[20] = `CIPHERTEXT_WIDTH'd11431889;
cipher_text[21] = `CIPHERTEXT_WIDTH'd12436186;
cipher_text[22] = `CIPHERTEXT_WIDTH'd4884439;
cipher_text[23] = `CIPHERTEXT_WIDTH'd12034802;
cipher_text[24] = `CIPHERTEXT_WIDTH'd605134;
cipher_text[25] = `CIPHERTEXT_WIDTH'd7252483;
cipher_text[26] = `CIPHERTEXT_WIDTH'd5544777;
cipher_text[27] = `CIPHERTEXT_WIDTH'd2132429;
cipher_text[28] = `CIPHERTEXT_WIDTH'd14207448;
cipher_text[29] = `CIPHERTEXT_WIDTH'd3427142;
cipher_text[30] = `CIPHERTEXT_WIDTH'd12814586;
cipher_text[31] = `CIPHERTEXT_WIDTH'd2282272;
cipher_text[32] = `CIPHERTEXT_WIDTH'd10458918;
cipher_text[33] = `CIPHERTEXT_WIDTH'd11087081;
cipher_text[34] = `CIPHERTEXT_WIDTH'd9384957;
cipher_text[35] = `CIPHERTEXT_WIDTH'd13802923;
cipher_text[36] = `CIPHERTEXT_WIDTH'd14314675;
cipher_text[37] = `CIPHERTEXT_WIDTH'd14616397;
cipher_text[38] = `CIPHERTEXT_WIDTH'd16379271;
cipher_text[39] = `CIPHERTEXT_WIDTH'd10427720;
cipher_text[40] = `CIPHERTEXT_WIDTH'd1014720;
cipher_text[41] = `CIPHERTEXT_WIDTH'd12583343;
cipher_text[42] = `CIPHERTEXT_WIDTH'd7993497;
cipher_text[43] = `CIPHERTEXT_WIDTH'd14460511;
cipher_text[44] = `CIPHERTEXT_WIDTH'd544346;
cipher_text[45] = `CIPHERTEXT_WIDTH'd8117013;
cipher_text[46] = `CIPHERTEXT_WIDTH'd4826204;
cipher_text[47] = `CIPHERTEXT_WIDTH'd16093233;
cipher_text[48] = `CIPHERTEXT_WIDTH'd6129358;
cipher_text[49] = `CIPHERTEXT_WIDTH'd9620921;
cipher_text[50] = `CIPHERTEXT_WIDTH'd13646236;
cipher_text[51] = `CIPHERTEXT_WIDTH'd3235218;
cipher_text[52] = `CIPHERTEXT_WIDTH'd1735224;
cipher_text[53] = `CIPHERTEXT_WIDTH'd109276;
cipher_text[54] = `CIPHERTEXT_WIDTH'd2489800;
cipher_text[55] = `CIPHERTEXT_WIDTH'd1849574;
cipher_text[56] = `CIPHERTEXT_WIDTH'd2315573;
cipher_text[57] = `CIPHERTEXT_WIDTH'd11071608;
cipher_text[58] = `CIPHERTEXT_WIDTH'd1252165;
cipher_text[59] = `CIPHERTEXT_WIDTH'd13185328;
cipher_text[60] = `CIPHERTEXT_WIDTH'd68417;
cipher_text[61] = `CIPHERTEXT_WIDTH'd3183599;
cipher_text[62] = `CIPHERTEXT_WIDTH'd15552599;
cipher_text[63] = `CIPHERTEXT_WIDTH'd15347029;
cipher_text[64] = `CIPHERTEXT_WIDTH'd12203675;
cipher_text[65] = `CIPHERTEXT_WIDTH'd2136663;
cipher_text[66] = `CIPHERTEXT_WIDTH'd12189268;
cipher_text[67] = `CIPHERTEXT_WIDTH'd7858238;
cipher_text[68] = `CIPHERTEXT_WIDTH'd5002646;
cipher_text[69] = `CIPHERTEXT_WIDTH'd6036590;
cipher_text[70] = `CIPHERTEXT_WIDTH'd1707794;
cipher_text[71] = `CIPHERTEXT_WIDTH'd12007582;
cipher_text[72] = `CIPHERTEXT_WIDTH'd14933659;
cipher_text[73] = `CIPHERTEXT_WIDTH'd8326192;
cipher_text[74] = `CIPHERTEXT_WIDTH'd6071656;
cipher_text[75] = `CIPHERTEXT_WIDTH'd15709017;
cipher_text[76] = `CIPHERTEXT_WIDTH'd9815848;
cipher_text[77] = `CIPHERTEXT_WIDTH'd6697436;
cipher_text[78] = `CIPHERTEXT_WIDTH'd188085;
cipher_text[79] = `CIPHERTEXT_WIDTH'd16236723;
cipher_text[80] = `CIPHERTEXT_WIDTH'd895125;
cipher_text[81] = `CIPHERTEXT_WIDTH'd6530206;
cipher_text[82] = `CIPHERTEXT_WIDTH'd11855117;
cipher_text[83] = `CIPHERTEXT_WIDTH'd11879029;
cipher_text[84] = `CIPHERTEXT_WIDTH'd5490857;
cipher_text[85] = `CIPHERTEXT_WIDTH'd11057928;
cipher_text[86] = `CIPHERTEXT_WIDTH'd7661666;
cipher_text[87] = `CIPHERTEXT_WIDTH'd8864449;
cipher_text[88] = `CIPHERTEXT_WIDTH'd1034932;
cipher_text[89] = `CIPHERTEXT_WIDTH'd5792880;
cipher_text[90] = `CIPHERTEXT_WIDTH'd6283655;
cipher_text[91] = `CIPHERTEXT_WIDTH'd12899309;
cipher_text[92] = `CIPHERTEXT_WIDTH'd4498754;
cipher_text[93] = `CIPHERTEXT_WIDTH'd13592626;
cipher_text[94] = `CIPHERTEXT_WIDTH'd13389174;
cipher_text[95] = `CIPHERTEXT_WIDTH'd10222781;
cipher_text[96] = `CIPHERTEXT_WIDTH'd8320536;
cipher_text[97] = `CIPHERTEXT_WIDTH'd6753823;
cipher_text[98] = `CIPHERTEXT_WIDTH'd11426289;
cipher_text[99] = `CIPHERTEXT_WIDTH'd1576985;
cipher_text[100] = `CIPHERTEXT_WIDTH'd1819706;
cipher_text[101] = `CIPHERTEXT_WIDTH'd6736242;
cipher_text[102] = `CIPHERTEXT_WIDTH'd5213699;
cipher_text[103] = `CIPHERTEXT_WIDTH'd7651620;
cipher_text[104] = `CIPHERTEXT_WIDTH'd1387171;
cipher_text[105] = `CIPHERTEXT_WIDTH'd13227674;
cipher_text[106] = `CIPHERTEXT_WIDTH'd11738951;
cipher_text[107] = `CIPHERTEXT_WIDTH'd7916216;
cipher_text[108] = `CIPHERTEXT_WIDTH'd3708782;
cipher_text[109] = `CIPHERTEXT_WIDTH'd567226;
cipher_text[110] = `CIPHERTEXT_WIDTH'd10011852;
cipher_text[111] = `CIPHERTEXT_WIDTH'd12791334;
cipher_text[112] = `CIPHERTEXT_WIDTH'd5541111;
cipher_text[113] = `CIPHERTEXT_WIDTH'd6783927;
cipher_text[114] = `CIPHERTEXT_WIDTH'd12214199;
cipher_text[115] = `CIPHERTEXT_WIDTH'd1388595;
cipher_text[116] = `CIPHERTEXT_WIDTH'd13587655;
cipher_text[117] = `CIPHERTEXT_WIDTH'd11669603;
cipher_text[118] = `CIPHERTEXT_WIDTH'd8287069;
cipher_text[119] = `CIPHERTEXT_WIDTH'd7142729;
cipher_text[120] = `CIPHERTEXT_WIDTH'd11367939;
cipher_text[121] = `CIPHERTEXT_WIDTH'd16333460;
cipher_text[122] = `CIPHERTEXT_WIDTH'd13191410;
cipher_text[123] = `CIPHERTEXT_WIDTH'd12374348;
cipher_text[124] = `CIPHERTEXT_WIDTH'd12245347;
cipher_text[125] = `CIPHERTEXT_WIDTH'd15936030;
cipher_text[126] = `CIPHERTEXT_WIDTH'd107215;
cipher_text[127] = `CIPHERTEXT_WIDTH'd787897;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 1;
cipher_text[0] = `CIPHERTEXT_WIDTH'd9865868;
cipher_text[1] = `CIPHERTEXT_WIDTH'd8932788;
cipher_text[2] = `CIPHERTEXT_WIDTH'd3588366;
cipher_text[3] = `CIPHERTEXT_WIDTH'd7923578;
cipher_text[4] = `CIPHERTEXT_WIDTH'd13393216;
cipher_text[5] = `CIPHERTEXT_WIDTH'd7523869;
cipher_text[6] = `CIPHERTEXT_WIDTH'd12548829;
cipher_text[7] = `CIPHERTEXT_WIDTH'd2634529;
cipher_text[8] = `CIPHERTEXT_WIDTH'd10205480;
cipher_text[9] = `CIPHERTEXT_WIDTH'd10027610;
cipher_text[10] = `CIPHERTEXT_WIDTH'd4688175;
cipher_text[11] = `CIPHERTEXT_WIDTH'd6612040;
cipher_text[12] = `CIPHERTEXT_WIDTH'd9385035;
cipher_text[13] = `CIPHERTEXT_WIDTH'd1116623;
cipher_text[14] = `CIPHERTEXT_WIDTH'd754361;
cipher_text[15] = `CIPHERTEXT_WIDTH'd5964592;
cipher_text[16] = `CIPHERTEXT_WIDTH'd4720989;
cipher_text[17] = `CIPHERTEXT_WIDTH'd1084887;
cipher_text[18] = `CIPHERTEXT_WIDTH'd11503306;
cipher_text[19] = `CIPHERTEXT_WIDTH'd10329481;
cipher_text[20] = `CIPHERTEXT_WIDTH'd12792553;
cipher_text[21] = `CIPHERTEXT_WIDTH'd3078936;
cipher_text[22] = `CIPHERTEXT_WIDTH'd13847651;
cipher_text[23] = `CIPHERTEXT_WIDTH'd12390560;
cipher_text[24] = `CIPHERTEXT_WIDTH'd11018654;
cipher_text[25] = `CIPHERTEXT_WIDTH'd7763659;
cipher_text[26] = `CIPHERTEXT_WIDTH'd9061711;
cipher_text[27] = `CIPHERTEXT_WIDTH'd10041338;
cipher_text[28] = `CIPHERTEXT_WIDTH'd16619535;
cipher_text[29] = `CIPHERTEXT_WIDTH'd5570667;
cipher_text[30] = `CIPHERTEXT_WIDTH'd3692402;
cipher_text[31] = `CIPHERTEXT_WIDTH'd15090947;
cipher_text[32] = `CIPHERTEXT_WIDTH'd340827;
cipher_text[33] = `CIPHERTEXT_WIDTH'd8294605;
cipher_text[34] = `CIPHERTEXT_WIDTH'd6208856;
cipher_text[35] = `CIPHERTEXT_WIDTH'd14303550;
cipher_text[36] = `CIPHERTEXT_WIDTH'd11762749;
cipher_text[37] = `CIPHERTEXT_WIDTH'd6192901;
cipher_text[38] = `CIPHERTEXT_WIDTH'd14784915;
cipher_text[39] = `CIPHERTEXT_WIDTH'd11009484;
cipher_text[40] = `CIPHERTEXT_WIDTH'd13976374;
cipher_text[41] = `CIPHERTEXT_WIDTH'd14299184;
cipher_text[42] = `CIPHERTEXT_WIDTH'd10389979;
cipher_text[43] = `CIPHERTEXT_WIDTH'd4697223;
cipher_text[44] = `CIPHERTEXT_WIDTH'd5870723;
cipher_text[45] = `CIPHERTEXT_WIDTH'd10430014;
cipher_text[46] = `CIPHERTEXT_WIDTH'd5806482;
cipher_text[47] = `CIPHERTEXT_WIDTH'd5387129;
cipher_text[48] = `CIPHERTEXT_WIDTH'd7410895;
cipher_text[49] = `CIPHERTEXT_WIDTH'd14124558;
cipher_text[50] = `CIPHERTEXT_WIDTH'd123349;
cipher_text[51] = `CIPHERTEXT_WIDTH'd15235460;
cipher_text[52] = `CIPHERTEXT_WIDTH'd5140136;
cipher_text[53] = `CIPHERTEXT_WIDTH'd12978688;
cipher_text[54] = `CIPHERTEXT_WIDTH'd4060529;
cipher_text[55] = `CIPHERTEXT_WIDTH'd2578706;
cipher_text[56] = `CIPHERTEXT_WIDTH'd6831350;
cipher_text[57] = `CIPHERTEXT_WIDTH'd10548151;
cipher_text[58] = `CIPHERTEXT_WIDTH'd12062771;
cipher_text[59] = `CIPHERTEXT_WIDTH'd6949453;
cipher_text[60] = `CIPHERTEXT_WIDTH'd6642264;
cipher_text[61] = `CIPHERTEXT_WIDTH'd9054259;
cipher_text[62] = `CIPHERTEXT_WIDTH'd9269070;
cipher_text[63] = `CIPHERTEXT_WIDTH'd9324384;
cipher_text[64] = `CIPHERTEXT_WIDTH'd187243;
cipher_text[65] = `CIPHERTEXT_WIDTH'd12012721;
cipher_text[66] = `CIPHERTEXT_WIDTH'd8001227;
cipher_text[67] = `CIPHERTEXT_WIDTH'd13027063;
cipher_text[68] = `CIPHERTEXT_WIDTH'd7982638;
cipher_text[69] = `CIPHERTEXT_WIDTH'd3545946;
cipher_text[70] = `CIPHERTEXT_WIDTH'd14396667;
cipher_text[71] = `CIPHERTEXT_WIDTH'd7999856;
cipher_text[72] = `CIPHERTEXT_WIDTH'd7679715;
cipher_text[73] = `CIPHERTEXT_WIDTH'd8632136;
cipher_text[74] = `CIPHERTEXT_WIDTH'd7012904;
cipher_text[75] = `CIPHERTEXT_WIDTH'd12139671;
cipher_text[76] = `CIPHERTEXT_WIDTH'd1772035;
cipher_text[77] = `CIPHERTEXT_WIDTH'd4797815;
cipher_text[78] = `CIPHERTEXT_WIDTH'd4634701;
cipher_text[79] = `CIPHERTEXT_WIDTH'd12237784;
cipher_text[80] = `CIPHERTEXT_WIDTH'd1754924;
cipher_text[81] = `CIPHERTEXT_WIDTH'd14729640;
cipher_text[82] = `CIPHERTEXT_WIDTH'd10660992;
cipher_text[83] = `CIPHERTEXT_WIDTH'd1413798;
cipher_text[84] = `CIPHERTEXT_WIDTH'd2127409;
cipher_text[85] = `CIPHERTEXT_WIDTH'd271150;
cipher_text[86] = `CIPHERTEXT_WIDTH'd14691086;
cipher_text[87] = `CIPHERTEXT_WIDTH'd7267069;
cipher_text[88] = `CIPHERTEXT_WIDTH'd14168743;
cipher_text[89] = `CIPHERTEXT_WIDTH'd2756859;
cipher_text[90] = `CIPHERTEXT_WIDTH'd10507909;
cipher_text[91] = `CIPHERTEXT_WIDTH'd1158605;
cipher_text[92] = `CIPHERTEXT_WIDTH'd2773851;
cipher_text[93] = `CIPHERTEXT_WIDTH'd12934378;
cipher_text[94] = `CIPHERTEXT_WIDTH'd5678103;
cipher_text[95] = `CIPHERTEXT_WIDTH'd2750165;
cipher_text[96] = `CIPHERTEXT_WIDTH'd14419799;
cipher_text[97] = `CIPHERTEXT_WIDTH'd8736394;
cipher_text[98] = `CIPHERTEXT_WIDTH'd16507934;
cipher_text[99] = `CIPHERTEXT_WIDTH'd1599732;
cipher_text[100] = `CIPHERTEXT_WIDTH'd5589789;
cipher_text[101] = `CIPHERTEXT_WIDTH'd2714260;
cipher_text[102] = `CIPHERTEXT_WIDTH'd5856304;
cipher_text[103] = `CIPHERTEXT_WIDTH'd7640440;
cipher_text[104] = `CIPHERTEXT_WIDTH'd13544276;
cipher_text[105] = `CIPHERTEXT_WIDTH'd13806186;
cipher_text[106] = `CIPHERTEXT_WIDTH'd15062071;
cipher_text[107] = `CIPHERTEXT_WIDTH'd9138667;
cipher_text[108] = `CIPHERTEXT_WIDTH'd14937982;
cipher_text[109] = `CIPHERTEXT_WIDTH'd14715247;
cipher_text[110] = `CIPHERTEXT_WIDTH'd8746041;
cipher_text[111] = `CIPHERTEXT_WIDTH'd12700632;
cipher_text[112] = `CIPHERTEXT_WIDTH'd13552955;
cipher_text[113] = `CIPHERTEXT_WIDTH'd4155876;
cipher_text[114] = `CIPHERTEXT_WIDTH'd16128585;
cipher_text[115] = `CIPHERTEXT_WIDTH'd14079732;
cipher_text[116] = `CIPHERTEXT_WIDTH'd9985688;
cipher_text[117] = `CIPHERTEXT_WIDTH'd5634802;
cipher_text[118] = `CIPHERTEXT_WIDTH'd9394681;
cipher_text[119] = `CIPHERTEXT_WIDTH'd11962686;
cipher_text[120] = `CIPHERTEXT_WIDTH'd11413530;
cipher_text[121] = `CIPHERTEXT_WIDTH'd15410613;
cipher_text[122] = `CIPHERTEXT_WIDTH'd10906515;
cipher_text[123] = `CIPHERTEXT_WIDTH'd7614069;
cipher_text[124] = `CIPHERTEXT_WIDTH'd13292621;
cipher_text[125] = `CIPHERTEXT_WIDTH'd16363252;
cipher_text[126] = `CIPHERTEXT_WIDTH'd16462111;
cipher_text[127] = `CIPHERTEXT_WIDTH'd15327814;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 2;
cipher_text[0] = `CIPHERTEXT_WIDTH'd1387670;
cipher_text[1] = `CIPHERTEXT_WIDTH'd3954895;
cipher_text[2] = `CIPHERTEXT_WIDTH'd15808792;
cipher_text[3] = `CIPHERTEXT_WIDTH'd13607405;
cipher_text[4] = `CIPHERTEXT_WIDTH'd16154900;
cipher_text[5] = `CIPHERTEXT_WIDTH'd2646115;
cipher_text[6] = `CIPHERTEXT_WIDTH'd16629226;
cipher_text[7] = `CIPHERTEXT_WIDTH'd13177082;
cipher_text[8] = `CIPHERTEXT_WIDTH'd8326980;
cipher_text[9] = `CIPHERTEXT_WIDTH'd5766200;
cipher_text[10] = `CIPHERTEXT_WIDTH'd225867;
cipher_text[11] = `CIPHERTEXT_WIDTH'd6655091;
cipher_text[12] = `CIPHERTEXT_WIDTH'd13958499;
cipher_text[13] = `CIPHERTEXT_WIDTH'd6147929;
cipher_text[14] = `CIPHERTEXT_WIDTH'd6413391;
cipher_text[15] = `CIPHERTEXT_WIDTH'd11801972;
cipher_text[16] = `CIPHERTEXT_WIDTH'd7529053;
cipher_text[17] = `CIPHERTEXT_WIDTH'd699814;
cipher_text[18] = `CIPHERTEXT_WIDTH'd6686461;
cipher_text[19] = `CIPHERTEXT_WIDTH'd11728974;
cipher_text[20] = `CIPHERTEXT_WIDTH'd11316959;
cipher_text[21] = `CIPHERTEXT_WIDTH'd1469787;
cipher_text[22] = `CIPHERTEXT_WIDTH'd4242735;
cipher_text[23] = `CIPHERTEXT_WIDTH'd1292947;
cipher_text[24] = `CIPHERTEXT_WIDTH'd15762412;
cipher_text[25] = `CIPHERTEXT_WIDTH'd2359930;
cipher_text[26] = `CIPHERTEXT_WIDTH'd16348537;
cipher_text[27] = `CIPHERTEXT_WIDTH'd3125765;
cipher_text[28] = `CIPHERTEXT_WIDTH'd13853217;
cipher_text[29] = `CIPHERTEXT_WIDTH'd7023750;
cipher_text[30] = `CIPHERTEXT_WIDTH'd12438748;
cipher_text[31] = `CIPHERTEXT_WIDTH'd1759331;
cipher_text[32] = `CIPHERTEXT_WIDTH'd4720805;
cipher_text[33] = `CIPHERTEXT_WIDTH'd2248658;
cipher_text[34] = `CIPHERTEXT_WIDTH'd3455108;
cipher_text[35] = `CIPHERTEXT_WIDTH'd16018236;
cipher_text[36] = `CIPHERTEXT_WIDTH'd2540011;
cipher_text[37] = `CIPHERTEXT_WIDTH'd9818189;
cipher_text[38] = `CIPHERTEXT_WIDTH'd3407169;
cipher_text[39] = `CIPHERTEXT_WIDTH'd8461847;
cipher_text[40] = `CIPHERTEXT_WIDTH'd3219667;
cipher_text[41] = `CIPHERTEXT_WIDTH'd15126085;
cipher_text[42] = `CIPHERTEXT_WIDTH'd14341081;
cipher_text[43] = `CIPHERTEXT_WIDTH'd2270075;
cipher_text[44] = `CIPHERTEXT_WIDTH'd8850877;
cipher_text[45] = `CIPHERTEXT_WIDTH'd5338038;
cipher_text[46] = `CIPHERTEXT_WIDTH'd568326;
cipher_text[47] = `CIPHERTEXT_WIDTH'd13669413;
cipher_text[48] = `CIPHERTEXT_WIDTH'd8788223;
cipher_text[49] = `CIPHERTEXT_WIDTH'd1217783;
cipher_text[50] = `CIPHERTEXT_WIDTH'd3679631;
cipher_text[51] = `CIPHERTEXT_WIDTH'd6116050;
cipher_text[52] = `CIPHERTEXT_WIDTH'd15356715;
cipher_text[53] = `CIPHERTEXT_WIDTH'd8388203;
cipher_text[54] = `CIPHERTEXT_WIDTH'd15450083;
cipher_text[55] = `CIPHERTEXT_WIDTH'd13377113;
cipher_text[56] = `CIPHERTEXT_WIDTH'd11752436;
cipher_text[57] = `CIPHERTEXT_WIDTH'd1924752;
cipher_text[58] = `CIPHERTEXT_WIDTH'd9507934;
cipher_text[59] = `CIPHERTEXT_WIDTH'd3682386;
cipher_text[60] = `CIPHERTEXT_WIDTH'd10778053;
cipher_text[61] = `CIPHERTEXT_WIDTH'd9480459;
cipher_text[62] = `CIPHERTEXT_WIDTH'd3726044;
cipher_text[63] = `CIPHERTEXT_WIDTH'd7324362;
cipher_text[64] = `CIPHERTEXT_WIDTH'd4434710;
cipher_text[65] = `CIPHERTEXT_WIDTH'd12110855;
cipher_text[66] = `CIPHERTEXT_WIDTH'd12474350;
cipher_text[67] = `CIPHERTEXT_WIDTH'd3476649;
cipher_text[68] = `CIPHERTEXT_WIDTH'd6930821;
cipher_text[69] = `CIPHERTEXT_WIDTH'd16774579;
cipher_text[70] = `CIPHERTEXT_WIDTH'd348642;
cipher_text[71] = `CIPHERTEXT_WIDTH'd14331415;
cipher_text[72] = `CIPHERTEXT_WIDTH'd9000315;
cipher_text[73] = `CIPHERTEXT_WIDTH'd12146297;
cipher_text[74] = `CIPHERTEXT_WIDTH'd3750795;
cipher_text[75] = `CIPHERTEXT_WIDTH'd11225611;
cipher_text[76] = `CIPHERTEXT_WIDTH'd8466458;
cipher_text[77] = `CIPHERTEXT_WIDTH'd2914574;
cipher_text[78] = `CIPHERTEXT_WIDTH'd243503;
cipher_text[79] = `CIPHERTEXT_WIDTH'd10639959;
cipher_text[80] = `CIPHERTEXT_WIDTH'd14598676;
cipher_text[81] = `CIPHERTEXT_WIDTH'd3515017;
cipher_text[82] = `CIPHERTEXT_WIDTH'd2886278;
cipher_text[83] = `CIPHERTEXT_WIDTH'd11259006;
cipher_text[84] = `CIPHERTEXT_WIDTH'd8826906;
cipher_text[85] = `CIPHERTEXT_WIDTH'd2006231;
cipher_text[86] = `CIPHERTEXT_WIDTH'd750727;
cipher_text[87] = `CIPHERTEXT_WIDTH'd12742386;
cipher_text[88] = `CIPHERTEXT_WIDTH'd12062851;
cipher_text[89] = `CIPHERTEXT_WIDTH'd14319674;
cipher_text[90] = `CIPHERTEXT_WIDTH'd15917958;
cipher_text[91] = `CIPHERTEXT_WIDTH'd12973852;
cipher_text[92] = `CIPHERTEXT_WIDTH'd15316311;
cipher_text[93] = `CIPHERTEXT_WIDTH'd7149739;
cipher_text[94] = `CIPHERTEXT_WIDTH'd13327516;
cipher_text[95] = `CIPHERTEXT_WIDTH'd14349133;
cipher_text[96] = `CIPHERTEXT_WIDTH'd15687225;
cipher_text[97] = `CIPHERTEXT_WIDTH'd3189323;
cipher_text[98] = `CIPHERTEXT_WIDTH'd15316804;
cipher_text[99] = `CIPHERTEXT_WIDTH'd6006656;
cipher_text[100] = `CIPHERTEXT_WIDTH'd26129;
cipher_text[101] = `CIPHERTEXT_WIDTH'd5262995;
cipher_text[102] = `CIPHERTEXT_WIDTH'd123764;
cipher_text[103] = `CIPHERTEXT_WIDTH'd6435607;
cipher_text[104] = `CIPHERTEXT_WIDTH'd1488270;
cipher_text[105] = `CIPHERTEXT_WIDTH'd13699372;
cipher_text[106] = `CIPHERTEXT_WIDTH'd16678271;
cipher_text[107] = `CIPHERTEXT_WIDTH'd4648510;
cipher_text[108] = `CIPHERTEXT_WIDTH'd15866854;
cipher_text[109] = `CIPHERTEXT_WIDTH'd14590858;
cipher_text[110] = `CIPHERTEXT_WIDTH'd15126500;
cipher_text[111] = `CIPHERTEXT_WIDTH'd7545884;
cipher_text[112] = `CIPHERTEXT_WIDTH'd8315322;
cipher_text[113] = `CIPHERTEXT_WIDTH'd13311672;
cipher_text[114] = `CIPHERTEXT_WIDTH'd10176983;
cipher_text[115] = `CIPHERTEXT_WIDTH'd4598564;
cipher_text[116] = `CIPHERTEXT_WIDTH'd16071498;
cipher_text[117] = `CIPHERTEXT_WIDTH'd77253;
cipher_text[118] = `CIPHERTEXT_WIDTH'd6504068;
cipher_text[119] = `CIPHERTEXT_WIDTH'd9397754;
cipher_text[120] = `CIPHERTEXT_WIDTH'd1879720;
cipher_text[121] = `CIPHERTEXT_WIDTH'd13110755;
cipher_text[122] = `CIPHERTEXT_WIDTH'd5476373;
cipher_text[123] = `CIPHERTEXT_WIDTH'd8544490;
cipher_text[124] = `CIPHERTEXT_WIDTH'd12337977;
cipher_text[125] = `CIPHERTEXT_WIDTH'd7966827;
cipher_text[126] = `CIPHERTEXT_WIDTH'd2169156;
cipher_text[127] = `CIPHERTEXT_WIDTH'd11472090;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 3;
cipher_text[0] = `CIPHERTEXT_WIDTH'd9007224;
cipher_text[1] = `CIPHERTEXT_WIDTH'd5415436;
cipher_text[2] = `CIPHERTEXT_WIDTH'd3895050;
cipher_text[3] = `CIPHERTEXT_WIDTH'd8930083;
cipher_text[4] = `CIPHERTEXT_WIDTH'd1688424;
cipher_text[5] = `CIPHERTEXT_WIDTH'd12150230;
cipher_text[6] = `CIPHERTEXT_WIDTH'd14908343;
cipher_text[7] = `CIPHERTEXT_WIDTH'd3178208;
cipher_text[8] = `CIPHERTEXT_WIDTH'd16400682;
cipher_text[9] = `CIPHERTEXT_WIDTH'd7191644;
cipher_text[10] = `CIPHERTEXT_WIDTH'd2786560;
cipher_text[11] = `CIPHERTEXT_WIDTH'd13716814;
cipher_text[12] = `CIPHERTEXT_WIDTH'd9152940;
cipher_text[13] = `CIPHERTEXT_WIDTH'd6973512;
cipher_text[14] = `CIPHERTEXT_WIDTH'd2772287;
cipher_text[15] = `CIPHERTEXT_WIDTH'd6390312;
cipher_text[16] = `CIPHERTEXT_WIDTH'd2800755;
cipher_text[17] = `CIPHERTEXT_WIDTH'd11955588;
cipher_text[18] = `CIPHERTEXT_WIDTH'd15808464;
cipher_text[19] = `CIPHERTEXT_WIDTH'd5646229;
cipher_text[20] = `CIPHERTEXT_WIDTH'd3801500;
cipher_text[21] = `CIPHERTEXT_WIDTH'd12896024;
cipher_text[22] = `CIPHERTEXT_WIDTH'd2051457;
cipher_text[23] = `CIPHERTEXT_WIDTH'd9210593;
cipher_text[24] = `CIPHERTEXT_WIDTH'd1220646;
cipher_text[25] = `CIPHERTEXT_WIDTH'd12330962;
cipher_text[26] = `CIPHERTEXT_WIDTH'd5413220;
cipher_text[27] = `CIPHERTEXT_WIDTH'd2231429;
cipher_text[28] = `CIPHERTEXT_WIDTH'd2806946;
cipher_text[29] = `CIPHERTEXT_WIDTH'd13966974;
cipher_text[30] = `CIPHERTEXT_WIDTH'd15865127;
cipher_text[31] = `CIPHERTEXT_WIDTH'd2798918;
cipher_text[32] = `CIPHERTEXT_WIDTH'd14602351;
cipher_text[33] = `CIPHERTEXT_WIDTH'd2429782;
cipher_text[34] = `CIPHERTEXT_WIDTH'd15481558;
cipher_text[35] = `CIPHERTEXT_WIDTH'd7367642;
cipher_text[36] = `CIPHERTEXT_WIDTH'd9275585;
cipher_text[37] = `CIPHERTEXT_WIDTH'd2779697;
cipher_text[38] = `CIPHERTEXT_WIDTH'd12355963;
cipher_text[39] = `CIPHERTEXT_WIDTH'd5451075;
cipher_text[40] = `CIPHERTEXT_WIDTH'd1988273;
cipher_text[41] = `CIPHERTEXT_WIDTH'd1773544;
cipher_text[42] = `CIPHERTEXT_WIDTH'd1264438;
cipher_text[43] = `CIPHERTEXT_WIDTH'd8312740;
cipher_text[44] = `CIPHERTEXT_WIDTH'd10023244;
cipher_text[45] = `CIPHERTEXT_WIDTH'd12748567;
cipher_text[46] = `CIPHERTEXT_WIDTH'd12260191;
cipher_text[47] = `CIPHERTEXT_WIDTH'd4067798;
cipher_text[48] = `CIPHERTEXT_WIDTH'd8875059;
cipher_text[49] = `CIPHERTEXT_WIDTH'd14952382;
cipher_text[50] = `CIPHERTEXT_WIDTH'd1174716;
cipher_text[51] = `CIPHERTEXT_WIDTH'd155849;
cipher_text[52] = `CIPHERTEXT_WIDTH'd7475013;
cipher_text[53] = `CIPHERTEXT_WIDTH'd9253169;
cipher_text[54] = `CIPHERTEXT_WIDTH'd15753522;
cipher_text[55] = `CIPHERTEXT_WIDTH'd9657691;
cipher_text[56] = `CIPHERTEXT_WIDTH'd7074337;
cipher_text[57] = `CIPHERTEXT_WIDTH'd1650603;
cipher_text[58] = `CIPHERTEXT_WIDTH'd6637692;
cipher_text[59] = `CIPHERTEXT_WIDTH'd4273589;
cipher_text[60] = `CIPHERTEXT_WIDTH'd9932580;
cipher_text[61] = `CIPHERTEXT_WIDTH'd2517258;
cipher_text[62] = `CIPHERTEXT_WIDTH'd12690287;
cipher_text[63] = `CIPHERTEXT_WIDTH'd13105015;
cipher_text[64] = `CIPHERTEXT_WIDTH'd3676685;
cipher_text[65] = `CIPHERTEXT_WIDTH'd5025324;
cipher_text[66] = `CIPHERTEXT_WIDTH'd16619523;
cipher_text[67] = `CIPHERTEXT_WIDTH'd12457053;
cipher_text[68] = `CIPHERTEXT_WIDTH'd479638;
cipher_text[69] = `CIPHERTEXT_WIDTH'd4429587;
cipher_text[70] = `CIPHERTEXT_WIDTH'd8749251;
cipher_text[71] = `CIPHERTEXT_WIDTH'd5412113;
cipher_text[72] = `CIPHERTEXT_WIDTH'd5128735;
cipher_text[73] = `CIPHERTEXT_WIDTH'd9682590;
cipher_text[74] = `CIPHERTEXT_WIDTH'd6229196;
cipher_text[75] = `CIPHERTEXT_WIDTH'd11010935;
cipher_text[76] = `CIPHERTEXT_WIDTH'd4994065;
cipher_text[77] = `CIPHERTEXT_WIDTH'd11466265;
cipher_text[78] = `CIPHERTEXT_WIDTH'd869;
cipher_text[79] = `CIPHERTEXT_WIDTH'd13444539;
cipher_text[80] = `CIPHERTEXT_WIDTH'd4384630;
cipher_text[81] = `CIPHERTEXT_WIDTH'd294543;
cipher_text[82] = `CIPHERTEXT_WIDTH'd290552;
cipher_text[83] = `CIPHERTEXT_WIDTH'd995465;
cipher_text[84] = `CIPHERTEXT_WIDTH'd2644886;
cipher_text[85] = `CIPHERTEXT_WIDTH'd13220984;
cipher_text[86] = `CIPHERTEXT_WIDTH'd4627745;
cipher_text[87] = `CIPHERTEXT_WIDTH'd859384;
cipher_text[88] = `CIPHERTEXT_WIDTH'd11140107;
cipher_text[89] = `CIPHERTEXT_WIDTH'd6818684;
cipher_text[90] = `CIPHERTEXT_WIDTH'd4135720;
cipher_text[91] = `CIPHERTEXT_WIDTH'd5687438;
cipher_text[92] = `CIPHERTEXT_WIDTH'd11165123;
cipher_text[93] = `CIPHERTEXT_WIDTH'd12820585;
cipher_text[94] = `CIPHERTEXT_WIDTH'd6876080;
cipher_text[95] = `CIPHERTEXT_WIDTH'd16117333;
cipher_text[96] = `CIPHERTEXT_WIDTH'd2820984;
cipher_text[97] = `CIPHERTEXT_WIDTH'd3729483;
cipher_text[98] = `CIPHERTEXT_WIDTH'd11204520;
cipher_text[99] = `CIPHERTEXT_WIDTH'd10830286;
cipher_text[100] = `CIPHERTEXT_WIDTH'd1640605;
cipher_text[101] = `CIPHERTEXT_WIDTH'd16493962;
cipher_text[102] = `CIPHERTEXT_WIDTH'd1696710;
cipher_text[103] = `CIPHERTEXT_WIDTH'd14236360;
cipher_text[104] = `CIPHERTEXT_WIDTH'd1859082;
cipher_text[105] = `CIPHERTEXT_WIDTH'd11977744;
cipher_text[106] = `CIPHERTEXT_WIDTH'd6630508;
cipher_text[107] = `CIPHERTEXT_WIDTH'd8414899;
cipher_text[108] = `CIPHERTEXT_WIDTH'd13677325;
cipher_text[109] = `CIPHERTEXT_WIDTH'd3227606;
cipher_text[110] = `CIPHERTEXT_WIDTH'd15278764;
cipher_text[111] = `CIPHERTEXT_WIDTH'd3420200;
cipher_text[112] = `CIPHERTEXT_WIDTH'd7361915;
cipher_text[113] = `CIPHERTEXT_WIDTH'd2924832;
cipher_text[114] = `CIPHERTEXT_WIDTH'd7397750;
cipher_text[115] = `CIPHERTEXT_WIDTH'd4467947;
cipher_text[116] = `CIPHERTEXT_WIDTH'd2243715;
cipher_text[117] = `CIPHERTEXT_WIDTH'd5246316;
cipher_text[118] = `CIPHERTEXT_WIDTH'd10433633;
cipher_text[119] = `CIPHERTEXT_WIDTH'd8993555;
cipher_text[120] = `CIPHERTEXT_WIDTH'd7856752;
cipher_text[121] = `CIPHERTEXT_WIDTH'd10339218;
cipher_text[122] = `CIPHERTEXT_WIDTH'd9956160;
cipher_text[123] = `CIPHERTEXT_WIDTH'd9554018;
cipher_text[124] = `CIPHERTEXT_WIDTH'd16657504;
cipher_text[125] = `CIPHERTEXT_WIDTH'd9160416;
cipher_text[126] = `CIPHERTEXT_WIDTH'd12114389;
cipher_text[127] = `CIPHERTEXT_WIDTH'd4135111;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 4;
cipher_text[0] = `CIPHERTEXT_WIDTH'd12114576;
cipher_text[1] = `CIPHERTEXT_WIDTH'd16446802;
cipher_text[2] = `CIPHERTEXT_WIDTH'd16161359;
cipher_text[3] = `CIPHERTEXT_WIDTH'd16343353;
cipher_text[4] = `CIPHERTEXT_WIDTH'd1681184;
cipher_text[5] = `CIPHERTEXT_WIDTH'd2210010;
cipher_text[6] = `CIPHERTEXT_WIDTH'd15318828;
cipher_text[7] = `CIPHERTEXT_WIDTH'd10430016;
cipher_text[8] = `CIPHERTEXT_WIDTH'd11233956;
cipher_text[9] = `CIPHERTEXT_WIDTH'd15202503;
cipher_text[10] = `CIPHERTEXT_WIDTH'd14928486;
cipher_text[11] = `CIPHERTEXT_WIDTH'd8434931;
cipher_text[12] = `CIPHERTEXT_WIDTH'd1379355;
cipher_text[13] = `CIPHERTEXT_WIDTH'd16142780;
cipher_text[14] = `CIPHERTEXT_WIDTH'd1850853;
cipher_text[15] = `CIPHERTEXT_WIDTH'd14235425;
cipher_text[16] = `CIPHERTEXT_WIDTH'd2826671;
cipher_text[17] = `CIPHERTEXT_WIDTH'd9794348;
cipher_text[18] = `CIPHERTEXT_WIDTH'd7234340;
cipher_text[19] = `CIPHERTEXT_WIDTH'd7033418;
cipher_text[20] = `CIPHERTEXT_WIDTH'd1797646;
cipher_text[21] = `CIPHERTEXT_WIDTH'd4882129;
cipher_text[22] = `CIPHERTEXT_WIDTH'd4694484;
cipher_text[23] = `CIPHERTEXT_WIDTH'd7139065;
cipher_text[24] = `CIPHERTEXT_WIDTH'd15994191;
cipher_text[25] = `CIPHERTEXT_WIDTH'd16402722;
cipher_text[26] = `CIPHERTEXT_WIDTH'd11066024;
cipher_text[27] = `CIPHERTEXT_WIDTH'd4215880;
cipher_text[28] = `CIPHERTEXT_WIDTH'd5296832;
cipher_text[29] = `CIPHERTEXT_WIDTH'd16406718;
cipher_text[30] = `CIPHERTEXT_WIDTH'd8296959;
cipher_text[31] = `CIPHERTEXT_WIDTH'd3505624;
cipher_text[32] = `CIPHERTEXT_WIDTH'd5091155;
cipher_text[33] = `CIPHERTEXT_WIDTH'd9276782;
cipher_text[34] = `CIPHERTEXT_WIDTH'd3659909;
cipher_text[35] = `CIPHERTEXT_WIDTH'd10556413;
cipher_text[36] = `CIPHERTEXT_WIDTH'd3664594;
cipher_text[37] = `CIPHERTEXT_WIDTH'd6200367;
cipher_text[38] = `CIPHERTEXT_WIDTH'd15496847;
cipher_text[39] = `CIPHERTEXT_WIDTH'd13452534;
cipher_text[40] = `CIPHERTEXT_WIDTH'd815698;
cipher_text[41] = `CIPHERTEXT_WIDTH'd3425235;
cipher_text[42] = `CIPHERTEXT_WIDTH'd14241723;
cipher_text[43] = `CIPHERTEXT_WIDTH'd10574796;
cipher_text[44] = `CIPHERTEXT_WIDTH'd14050545;
cipher_text[45] = `CIPHERTEXT_WIDTH'd2993443;
cipher_text[46] = `CIPHERTEXT_WIDTH'd11001874;
cipher_text[47] = `CIPHERTEXT_WIDTH'd283360;
cipher_text[48] = `CIPHERTEXT_WIDTH'd11166048;
cipher_text[49] = `CIPHERTEXT_WIDTH'd12955214;
cipher_text[50] = `CIPHERTEXT_WIDTH'd11552325;
cipher_text[51] = `CIPHERTEXT_WIDTH'd7836100;
cipher_text[52] = `CIPHERTEXT_WIDTH'd248151;
cipher_text[53] = `CIPHERTEXT_WIDTH'd7465535;
cipher_text[54] = `CIPHERTEXT_WIDTH'd7120769;
cipher_text[55] = `CIPHERTEXT_WIDTH'd13447523;
cipher_text[56] = `CIPHERTEXT_WIDTH'd6783802;
cipher_text[57] = `CIPHERTEXT_WIDTH'd14517514;
cipher_text[58] = `CIPHERTEXT_WIDTH'd6719110;
cipher_text[59] = `CIPHERTEXT_WIDTH'd2291368;
cipher_text[60] = `CIPHERTEXT_WIDTH'd13451545;
cipher_text[61] = `CIPHERTEXT_WIDTH'd12464917;
cipher_text[62] = `CIPHERTEXT_WIDTH'd6184591;
cipher_text[63] = `CIPHERTEXT_WIDTH'd12084071;
cipher_text[64] = `CIPHERTEXT_WIDTH'd16734401;
cipher_text[65] = `CIPHERTEXT_WIDTH'd1245237;
cipher_text[66] = `CIPHERTEXT_WIDTH'd5288848;
cipher_text[67] = `CIPHERTEXT_WIDTH'd15617581;
cipher_text[68] = `CIPHERTEXT_WIDTH'd13625669;
cipher_text[69] = `CIPHERTEXT_WIDTH'd11038626;
cipher_text[70] = `CIPHERTEXT_WIDTH'd16589425;
cipher_text[71] = `CIPHERTEXT_WIDTH'd7323319;
cipher_text[72] = `CIPHERTEXT_WIDTH'd14564737;
cipher_text[73] = `CIPHERTEXT_WIDTH'd11470805;
cipher_text[74] = `CIPHERTEXT_WIDTH'd11546366;
cipher_text[75] = `CIPHERTEXT_WIDTH'd11270836;
cipher_text[76] = `CIPHERTEXT_WIDTH'd5906082;
cipher_text[77] = `CIPHERTEXT_WIDTH'd513422;
cipher_text[78] = `CIPHERTEXT_WIDTH'd13209630;
cipher_text[79] = `CIPHERTEXT_WIDTH'd8098296;
cipher_text[80] = `CIPHERTEXT_WIDTH'd4075395;
cipher_text[81] = `CIPHERTEXT_WIDTH'd9925988;
cipher_text[82] = `CIPHERTEXT_WIDTH'd6385729;
cipher_text[83] = `CIPHERTEXT_WIDTH'd15573647;
cipher_text[84] = `CIPHERTEXT_WIDTH'd13416079;
cipher_text[85] = `CIPHERTEXT_WIDTH'd6799345;
cipher_text[86] = `CIPHERTEXT_WIDTH'd1510353;
cipher_text[87] = `CIPHERTEXT_WIDTH'd10231344;
cipher_text[88] = `CIPHERTEXT_WIDTH'd4324555;
cipher_text[89] = `CIPHERTEXT_WIDTH'd11426160;
cipher_text[90] = `CIPHERTEXT_WIDTH'd13996703;
cipher_text[91] = `CIPHERTEXT_WIDTH'd9578453;
cipher_text[92] = `CIPHERTEXT_WIDTH'd9482090;
cipher_text[93] = `CIPHERTEXT_WIDTH'd11343590;
cipher_text[94] = `CIPHERTEXT_WIDTH'd7576584;
cipher_text[95] = `CIPHERTEXT_WIDTH'd4778540;
cipher_text[96] = `CIPHERTEXT_WIDTH'd13311471;
cipher_text[97] = `CIPHERTEXT_WIDTH'd11556818;
cipher_text[98] = `CIPHERTEXT_WIDTH'd617576;
cipher_text[99] = `CIPHERTEXT_WIDTH'd4292688;
cipher_text[100] = `CIPHERTEXT_WIDTH'd3780458;
cipher_text[101] = `CIPHERTEXT_WIDTH'd14926527;
cipher_text[102] = `CIPHERTEXT_WIDTH'd16560650;
cipher_text[103] = `CIPHERTEXT_WIDTH'd3900709;
cipher_text[104] = `CIPHERTEXT_WIDTH'd16421798;
cipher_text[105] = `CIPHERTEXT_WIDTH'd9202286;
cipher_text[106] = `CIPHERTEXT_WIDTH'd16535260;
cipher_text[107] = `CIPHERTEXT_WIDTH'd3367504;
cipher_text[108] = `CIPHERTEXT_WIDTH'd13954447;
cipher_text[109] = `CIPHERTEXT_WIDTH'd13489183;
cipher_text[110] = `CIPHERTEXT_WIDTH'd9842803;
cipher_text[111] = `CIPHERTEXT_WIDTH'd605092;
cipher_text[112] = `CIPHERTEXT_WIDTH'd4968683;
cipher_text[113] = `CIPHERTEXT_WIDTH'd9402051;
cipher_text[114] = `CIPHERTEXT_WIDTH'd3051301;
cipher_text[115] = `CIPHERTEXT_WIDTH'd4148290;
cipher_text[116] = `CIPHERTEXT_WIDTH'd13447223;
cipher_text[117] = `CIPHERTEXT_WIDTH'd10146490;
cipher_text[118] = `CIPHERTEXT_WIDTH'd12998368;
cipher_text[119] = `CIPHERTEXT_WIDTH'd5331508;
cipher_text[120] = `CIPHERTEXT_WIDTH'd1392719;
cipher_text[121] = `CIPHERTEXT_WIDTH'd13698562;
cipher_text[122] = `CIPHERTEXT_WIDTH'd11610408;
cipher_text[123] = `CIPHERTEXT_WIDTH'd1886777;
cipher_text[124] = `CIPHERTEXT_WIDTH'd9935972;
cipher_text[125] = `CIPHERTEXT_WIDTH'd13178009;
cipher_text[126] = `CIPHERTEXT_WIDTH'd10015174;
cipher_text[127] = `CIPHERTEXT_WIDTH'd6564522;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 5;
cipher_text[0] = `CIPHERTEXT_WIDTH'd2920125;
cipher_text[1] = `CIPHERTEXT_WIDTH'd11363760;
cipher_text[2] = `CIPHERTEXT_WIDTH'd11558002;
cipher_text[3] = `CIPHERTEXT_WIDTH'd15918852;
cipher_text[4] = `CIPHERTEXT_WIDTH'd15905455;
cipher_text[5] = `CIPHERTEXT_WIDTH'd3842896;
cipher_text[6] = `CIPHERTEXT_WIDTH'd15009775;
cipher_text[7] = `CIPHERTEXT_WIDTH'd14692941;
cipher_text[8] = `CIPHERTEXT_WIDTH'd6468059;
cipher_text[9] = `CIPHERTEXT_WIDTH'd11120027;
cipher_text[10] = `CIPHERTEXT_WIDTH'd14485001;
cipher_text[11] = `CIPHERTEXT_WIDTH'd4430418;
cipher_text[12] = `CIPHERTEXT_WIDTH'd16112832;
cipher_text[13] = `CIPHERTEXT_WIDTH'd16383674;
cipher_text[14] = `CIPHERTEXT_WIDTH'd16385741;
cipher_text[15] = `CIPHERTEXT_WIDTH'd8669373;
cipher_text[16] = `CIPHERTEXT_WIDTH'd6263727;
cipher_text[17] = `CIPHERTEXT_WIDTH'd2828788;
cipher_text[18] = `CIPHERTEXT_WIDTH'd15674059;
cipher_text[19] = `CIPHERTEXT_WIDTH'd14455084;
cipher_text[20] = `CIPHERTEXT_WIDTH'd12399691;
cipher_text[21] = `CIPHERTEXT_WIDTH'd11325865;
cipher_text[22] = `CIPHERTEXT_WIDTH'd14697970;
cipher_text[23] = `CIPHERTEXT_WIDTH'd8221356;
cipher_text[24] = `CIPHERTEXT_WIDTH'd9544527;
cipher_text[25] = `CIPHERTEXT_WIDTH'd15455997;
cipher_text[26] = `CIPHERTEXT_WIDTH'd7285951;
cipher_text[27] = `CIPHERTEXT_WIDTH'd359404;
cipher_text[28] = `CIPHERTEXT_WIDTH'd7812388;
cipher_text[29] = `CIPHERTEXT_WIDTH'd6303639;
cipher_text[30] = `CIPHERTEXT_WIDTH'd6790125;
cipher_text[31] = `CIPHERTEXT_WIDTH'd3594583;
cipher_text[32] = `CIPHERTEXT_WIDTH'd3140963;
cipher_text[33] = `CIPHERTEXT_WIDTH'd11606581;
cipher_text[34] = `CIPHERTEXT_WIDTH'd11358949;
cipher_text[35] = `CIPHERTEXT_WIDTH'd14385631;
cipher_text[36] = `CIPHERTEXT_WIDTH'd13767140;
cipher_text[37] = `CIPHERTEXT_WIDTH'd277682;
cipher_text[38] = `CIPHERTEXT_WIDTH'd15375474;
cipher_text[39] = `CIPHERTEXT_WIDTH'd6391491;
cipher_text[40] = `CIPHERTEXT_WIDTH'd8210837;
cipher_text[41] = `CIPHERTEXT_WIDTH'd4135416;
cipher_text[42] = `CIPHERTEXT_WIDTH'd8822365;
cipher_text[43] = `CIPHERTEXT_WIDTH'd4237027;
cipher_text[44] = `CIPHERTEXT_WIDTH'd13607410;
cipher_text[45] = `CIPHERTEXT_WIDTH'd8282784;
cipher_text[46] = `CIPHERTEXT_WIDTH'd13261567;
cipher_text[47] = `CIPHERTEXT_WIDTH'd114293;
cipher_text[48] = `CIPHERTEXT_WIDTH'd8497474;
cipher_text[49] = `CIPHERTEXT_WIDTH'd4687659;
cipher_text[50] = `CIPHERTEXT_WIDTH'd5011351;
cipher_text[51] = `CIPHERTEXT_WIDTH'd16281967;
cipher_text[52] = `CIPHERTEXT_WIDTH'd7366012;
cipher_text[53] = `CIPHERTEXT_WIDTH'd13804702;
cipher_text[54] = `CIPHERTEXT_WIDTH'd10212001;
cipher_text[55] = `CIPHERTEXT_WIDTH'd5801894;
cipher_text[56] = `CIPHERTEXT_WIDTH'd244121;
cipher_text[57] = `CIPHERTEXT_WIDTH'd16078276;
cipher_text[58] = `CIPHERTEXT_WIDTH'd10256510;
cipher_text[59] = `CIPHERTEXT_WIDTH'd962118;
cipher_text[60] = `CIPHERTEXT_WIDTH'd8523623;
cipher_text[61] = `CIPHERTEXT_WIDTH'd930151;
cipher_text[62] = `CIPHERTEXT_WIDTH'd9952066;
cipher_text[63] = `CIPHERTEXT_WIDTH'd12638835;
cipher_text[64] = `CIPHERTEXT_WIDTH'd1108777;
cipher_text[65] = `CIPHERTEXT_WIDTH'd4123503;
cipher_text[66] = `CIPHERTEXT_WIDTH'd10382923;
cipher_text[67] = `CIPHERTEXT_WIDTH'd2034304;
cipher_text[68] = `CIPHERTEXT_WIDTH'd4324409;
cipher_text[69] = `CIPHERTEXT_WIDTH'd9453549;
cipher_text[70] = `CIPHERTEXT_WIDTH'd239988;
cipher_text[71] = `CIPHERTEXT_WIDTH'd15007630;
cipher_text[72] = `CIPHERTEXT_WIDTH'd5779559;
cipher_text[73] = `CIPHERTEXT_WIDTH'd2455974;
cipher_text[74] = `CIPHERTEXT_WIDTH'd15666816;
cipher_text[75] = `CIPHERTEXT_WIDTH'd816591;
cipher_text[76] = `CIPHERTEXT_WIDTH'd7202619;
cipher_text[77] = `CIPHERTEXT_WIDTH'd6307635;
cipher_text[78] = `CIPHERTEXT_WIDTH'd6653501;
cipher_text[79] = `CIPHERTEXT_WIDTH'd4712365;
cipher_text[80] = `CIPHERTEXT_WIDTH'd13494807;
cipher_text[81] = `CIPHERTEXT_WIDTH'd16598493;
cipher_text[82] = `CIPHERTEXT_WIDTH'd6496475;
cipher_text[83] = `CIPHERTEXT_WIDTH'd5442865;
cipher_text[84] = `CIPHERTEXT_WIDTH'd1923669;
cipher_text[85] = `CIPHERTEXT_WIDTH'd11680570;
cipher_text[86] = `CIPHERTEXT_WIDTH'd13278958;
cipher_text[87] = `CIPHERTEXT_WIDTH'd8331796;
cipher_text[88] = `CIPHERTEXT_WIDTH'd1622247;
cipher_text[89] = `CIPHERTEXT_WIDTH'd16281731;
cipher_text[90] = `CIPHERTEXT_WIDTH'd823864;
cipher_text[91] = `CIPHERTEXT_WIDTH'd312525;
cipher_text[92] = `CIPHERTEXT_WIDTH'd8727566;
cipher_text[93] = `CIPHERTEXT_WIDTH'd4272207;
cipher_text[94] = `CIPHERTEXT_WIDTH'd14453931;
cipher_text[95] = `CIPHERTEXT_WIDTH'd11581300;
cipher_text[96] = `CIPHERTEXT_WIDTH'd10934704;
cipher_text[97] = `CIPHERTEXT_WIDTH'd108926;
cipher_text[98] = `CIPHERTEXT_WIDTH'd13433673;
cipher_text[99] = `CIPHERTEXT_WIDTH'd5622559;
cipher_text[100] = `CIPHERTEXT_WIDTH'd14107501;
cipher_text[101] = `CIPHERTEXT_WIDTH'd8195126;
cipher_text[102] = `CIPHERTEXT_WIDTH'd13963716;
cipher_text[103] = `CIPHERTEXT_WIDTH'd8690729;
cipher_text[104] = `CIPHERTEXT_WIDTH'd9071134;
cipher_text[105] = `CIPHERTEXT_WIDTH'd10492042;
cipher_text[106] = `CIPHERTEXT_WIDTH'd14187797;
cipher_text[107] = `CIPHERTEXT_WIDTH'd16477363;
cipher_text[108] = `CIPHERTEXT_WIDTH'd6373527;
cipher_text[109] = `CIPHERTEXT_WIDTH'd271008;
cipher_text[110] = `CIPHERTEXT_WIDTH'd15792911;
cipher_text[111] = `CIPHERTEXT_WIDTH'd1128233;
cipher_text[112] = `CIPHERTEXT_WIDTH'd8652022;
cipher_text[113] = `CIPHERTEXT_WIDTH'd14529637;
cipher_text[114] = `CIPHERTEXT_WIDTH'd2613958;
cipher_text[115] = `CIPHERTEXT_WIDTH'd12481449;
cipher_text[116] = `CIPHERTEXT_WIDTH'd16718472;
cipher_text[117] = `CIPHERTEXT_WIDTH'd3923029;
cipher_text[118] = `CIPHERTEXT_WIDTH'd834481;
cipher_text[119] = `CIPHERTEXT_WIDTH'd1998770;
cipher_text[120] = `CIPHERTEXT_WIDTH'd15971156;
cipher_text[121] = `CIPHERTEXT_WIDTH'd12952244;
cipher_text[122] = `CIPHERTEXT_WIDTH'd13960327;
cipher_text[123] = `CIPHERTEXT_WIDTH'd1450716;
cipher_text[124] = `CIPHERTEXT_WIDTH'd16771396;
cipher_text[125] = `CIPHERTEXT_WIDTH'd4695715;
cipher_text[126] = `CIPHERTEXT_WIDTH'd1727154;
cipher_text[127] = `CIPHERTEXT_WIDTH'd1513968;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 6;
cipher_text[0] = `CIPHERTEXT_WIDTH'd3420591;
cipher_text[1] = `CIPHERTEXT_WIDTH'd5585276;
cipher_text[2] = `CIPHERTEXT_WIDTH'd6066620;
cipher_text[3] = `CIPHERTEXT_WIDTH'd1823398;
cipher_text[4] = `CIPHERTEXT_WIDTH'd1961788;
cipher_text[5] = `CIPHERTEXT_WIDTH'd8576972;
cipher_text[6] = `CIPHERTEXT_WIDTH'd5302829;
cipher_text[7] = `CIPHERTEXT_WIDTH'd8673668;
cipher_text[8] = `CIPHERTEXT_WIDTH'd6656829;
cipher_text[9] = `CIPHERTEXT_WIDTH'd10506277;
cipher_text[10] = `CIPHERTEXT_WIDTH'd11656608;
cipher_text[11] = `CIPHERTEXT_WIDTH'd9735112;
cipher_text[12] = `CIPHERTEXT_WIDTH'd4665254;
cipher_text[13] = `CIPHERTEXT_WIDTH'd16281113;
cipher_text[14] = `CIPHERTEXT_WIDTH'd4462845;
cipher_text[15] = `CIPHERTEXT_WIDTH'd5141603;
cipher_text[16] = `CIPHERTEXT_WIDTH'd14113975;
cipher_text[17] = `CIPHERTEXT_WIDTH'd6966566;
cipher_text[18] = `CIPHERTEXT_WIDTH'd14836754;
cipher_text[19] = `CIPHERTEXT_WIDTH'd2584614;
cipher_text[20] = `CIPHERTEXT_WIDTH'd827756;
cipher_text[21] = `CIPHERTEXT_WIDTH'd8645688;
cipher_text[22] = `CIPHERTEXT_WIDTH'd15744915;
cipher_text[23] = `CIPHERTEXT_WIDTH'd9002656;
cipher_text[24] = `CIPHERTEXT_WIDTH'd16348113;
cipher_text[25] = `CIPHERTEXT_WIDTH'd12377516;
cipher_text[26] = `CIPHERTEXT_WIDTH'd422345;
cipher_text[27] = `CIPHERTEXT_WIDTH'd12566663;
cipher_text[28] = `CIPHERTEXT_WIDTH'd10536752;
cipher_text[29] = `CIPHERTEXT_WIDTH'd13059259;
cipher_text[30] = `CIPHERTEXT_WIDTH'd1427408;
cipher_text[31] = `CIPHERTEXT_WIDTH'd5175449;
cipher_text[32] = `CIPHERTEXT_WIDTH'd14560183;
cipher_text[33] = `CIPHERTEXT_WIDTH'd8688810;
cipher_text[34] = `CIPHERTEXT_WIDTH'd7160765;
cipher_text[35] = `CIPHERTEXT_WIDTH'd7175305;
cipher_text[36] = `CIPHERTEXT_WIDTH'd9369623;
cipher_text[37] = `CIPHERTEXT_WIDTH'd13019542;
cipher_text[38] = `CIPHERTEXT_WIDTH'd14471354;
cipher_text[39] = `CIPHERTEXT_WIDTH'd6087830;
cipher_text[40] = `CIPHERTEXT_WIDTH'd6840733;
cipher_text[41] = `CIPHERTEXT_WIDTH'd7016858;
cipher_text[42] = `CIPHERTEXT_WIDTH'd9483474;
cipher_text[43] = `CIPHERTEXT_WIDTH'd4549880;
cipher_text[44] = `CIPHERTEXT_WIDTH'd10240691;
cipher_text[45] = `CIPHERTEXT_WIDTH'd4168113;
cipher_text[46] = `CIPHERTEXT_WIDTH'd2572658;
cipher_text[47] = `CIPHERTEXT_WIDTH'd8413636;
cipher_text[48] = `CIPHERTEXT_WIDTH'd11153631;
cipher_text[49] = `CIPHERTEXT_WIDTH'd8891073;
cipher_text[50] = `CIPHERTEXT_WIDTH'd4957154;
cipher_text[51] = `CIPHERTEXT_WIDTH'd4197559;
cipher_text[52] = `CIPHERTEXT_WIDTH'd10566608;
cipher_text[53] = `CIPHERTEXT_WIDTH'd4704506;
cipher_text[54] = `CIPHERTEXT_WIDTH'd204406;
cipher_text[55] = `CIPHERTEXT_WIDTH'd3109384;
cipher_text[56] = `CIPHERTEXT_WIDTH'd10138895;
cipher_text[57] = `CIPHERTEXT_WIDTH'd8745994;
cipher_text[58] = `CIPHERTEXT_WIDTH'd2951205;
cipher_text[59] = `CIPHERTEXT_WIDTH'd6599418;
cipher_text[60] = `CIPHERTEXT_WIDTH'd11532996;
cipher_text[61] = `CIPHERTEXT_WIDTH'd11943111;
cipher_text[62] = `CIPHERTEXT_WIDTH'd4973394;
cipher_text[63] = `CIPHERTEXT_WIDTH'd8115503;
cipher_text[64] = `CIPHERTEXT_WIDTH'd16564686;
cipher_text[65] = `CIPHERTEXT_WIDTH'd16518500;
cipher_text[66] = `CIPHERTEXT_WIDTH'd7260661;
cipher_text[67] = `CIPHERTEXT_WIDTH'd11245491;
cipher_text[68] = `CIPHERTEXT_WIDTH'd147667;
cipher_text[69] = `CIPHERTEXT_WIDTH'd7592846;
cipher_text[70] = `CIPHERTEXT_WIDTH'd47511;
cipher_text[71] = `CIPHERTEXT_WIDTH'd16298839;
cipher_text[72] = `CIPHERTEXT_WIDTH'd3318205;
cipher_text[73] = `CIPHERTEXT_WIDTH'd12259941;
cipher_text[74] = `CIPHERTEXT_WIDTH'd1845768;
cipher_text[75] = `CIPHERTEXT_WIDTH'd16335086;
cipher_text[76] = `CIPHERTEXT_WIDTH'd108758;
cipher_text[77] = `CIPHERTEXT_WIDTH'd326559;
cipher_text[78] = `CIPHERTEXT_WIDTH'd11353981;
cipher_text[79] = `CIPHERTEXT_WIDTH'd13838895;
cipher_text[80] = `CIPHERTEXT_WIDTH'd7172045;
cipher_text[81] = `CIPHERTEXT_WIDTH'd3552408;
cipher_text[82] = `CIPHERTEXT_WIDTH'd4475460;
cipher_text[83] = `CIPHERTEXT_WIDTH'd1846992;
cipher_text[84] = `CIPHERTEXT_WIDTH'd14010;
cipher_text[85] = `CIPHERTEXT_WIDTH'd1470178;
cipher_text[86] = `CIPHERTEXT_WIDTH'd15257722;
cipher_text[87] = `CIPHERTEXT_WIDTH'd13017227;
cipher_text[88] = `CIPHERTEXT_WIDTH'd2986912;
cipher_text[89] = `CIPHERTEXT_WIDTH'd1639813;
cipher_text[90] = `CIPHERTEXT_WIDTH'd5080346;
cipher_text[91] = `CIPHERTEXT_WIDTH'd6841524;
cipher_text[92] = `CIPHERTEXT_WIDTH'd5024118;
cipher_text[93] = `CIPHERTEXT_WIDTH'd12410121;
cipher_text[94] = `CIPHERTEXT_WIDTH'd15133406;
cipher_text[95] = `CIPHERTEXT_WIDTH'd13712372;
cipher_text[96] = `CIPHERTEXT_WIDTH'd10766947;
cipher_text[97] = `CIPHERTEXT_WIDTH'd14754029;
cipher_text[98] = `CIPHERTEXT_WIDTH'd9530128;
cipher_text[99] = `CIPHERTEXT_WIDTH'd9675475;
cipher_text[100] = `CIPHERTEXT_WIDTH'd3859727;
cipher_text[101] = `CIPHERTEXT_WIDTH'd12371614;
cipher_text[102] = `CIPHERTEXT_WIDTH'd1200140;
cipher_text[103] = `CIPHERTEXT_WIDTH'd2552621;
cipher_text[104] = `CIPHERTEXT_WIDTH'd12072296;
cipher_text[105] = `CIPHERTEXT_WIDTH'd4857315;
cipher_text[106] = `CIPHERTEXT_WIDTH'd11898875;
cipher_text[107] = `CIPHERTEXT_WIDTH'd3291794;
cipher_text[108] = `CIPHERTEXT_WIDTH'd4338288;
cipher_text[109] = `CIPHERTEXT_WIDTH'd5745610;
cipher_text[110] = `CIPHERTEXT_WIDTH'd4282012;
cipher_text[111] = `CIPHERTEXT_WIDTH'd9623292;
cipher_text[112] = `CIPHERTEXT_WIDTH'd2761305;
cipher_text[113] = `CIPHERTEXT_WIDTH'd1280800;
cipher_text[114] = `CIPHERTEXT_WIDTH'd4328287;
cipher_text[115] = `CIPHERTEXT_WIDTH'd13090593;
cipher_text[116] = `CIPHERTEXT_WIDTH'd7864479;
cipher_text[117] = `CIPHERTEXT_WIDTH'd10900617;
cipher_text[118] = `CIPHERTEXT_WIDTH'd10102455;
cipher_text[119] = `CIPHERTEXT_WIDTH'd8038524;
cipher_text[120] = `CIPHERTEXT_WIDTH'd4335781;
cipher_text[121] = `CIPHERTEXT_WIDTH'd4637887;
cipher_text[122] = `CIPHERTEXT_WIDTH'd7243424;
cipher_text[123] = `CIPHERTEXT_WIDTH'd12681010;
cipher_text[124] = `CIPHERTEXT_WIDTH'd10139096;
cipher_text[125] = `CIPHERTEXT_WIDTH'd115563;
cipher_text[126] = `CIPHERTEXT_WIDTH'd4381481;
cipher_text[127] = `CIPHERTEXT_WIDTH'd14385497;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 7;
cipher_text[0] = `CIPHERTEXT_WIDTH'd6454528;
cipher_text[1] = `CIPHERTEXT_WIDTH'd4355351;
cipher_text[2] = `CIPHERTEXT_WIDTH'd9775875;
cipher_text[3] = `CIPHERTEXT_WIDTH'd8125601;
cipher_text[4] = `CIPHERTEXT_WIDTH'd3064958;
cipher_text[5] = `CIPHERTEXT_WIDTH'd13286738;
cipher_text[6] = `CIPHERTEXT_WIDTH'd10601601;
cipher_text[7] = `CIPHERTEXT_WIDTH'd4071296;
cipher_text[8] = `CIPHERTEXT_WIDTH'd16231232;
cipher_text[9] = `CIPHERTEXT_WIDTH'd8787666;
cipher_text[10] = `CIPHERTEXT_WIDTH'd3072473;
cipher_text[11] = `CIPHERTEXT_WIDTH'd11653911;
cipher_text[12] = `CIPHERTEXT_WIDTH'd8553738;
cipher_text[13] = `CIPHERTEXT_WIDTH'd14679574;
cipher_text[14] = `CIPHERTEXT_WIDTH'd14726993;
cipher_text[15] = `CIPHERTEXT_WIDTH'd6628054;
cipher_text[16] = `CIPHERTEXT_WIDTH'd10321370;
cipher_text[17] = `CIPHERTEXT_WIDTH'd7632486;
cipher_text[18] = `CIPHERTEXT_WIDTH'd7635017;
cipher_text[19] = `CIPHERTEXT_WIDTH'd7758444;
cipher_text[20] = `CIPHERTEXT_WIDTH'd1660436;
cipher_text[21] = `CIPHERTEXT_WIDTH'd13255263;
cipher_text[22] = `CIPHERTEXT_WIDTH'd1637217;
cipher_text[23] = `CIPHERTEXT_WIDTH'd5357963;
cipher_text[24] = `CIPHERTEXT_WIDTH'd13610241;
cipher_text[25] = `CIPHERTEXT_WIDTH'd11349320;
cipher_text[26] = `CIPHERTEXT_WIDTH'd13678685;
cipher_text[27] = `CIPHERTEXT_WIDTH'd2313091;
cipher_text[28] = `CIPHERTEXT_WIDTH'd5084877;
cipher_text[29] = `CIPHERTEXT_WIDTH'd13905610;
cipher_text[30] = `CIPHERTEXT_WIDTH'd2725165;
cipher_text[31] = `CIPHERTEXT_WIDTH'd16191161;
cipher_text[32] = `CIPHERTEXT_WIDTH'd5450706;
cipher_text[33] = `CIPHERTEXT_WIDTH'd10510093;
cipher_text[34] = `CIPHERTEXT_WIDTH'd360069;
cipher_text[35] = `CIPHERTEXT_WIDTH'd15268004;
cipher_text[36] = `CIPHERTEXT_WIDTH'd9607656;
cipher_text[37] = `CIPHERTEXT_WIDTH'd12042100;
cipher_text[38] = `CIPHERTEXT_WIDTH'd7684779;
cipher_text[39] = `CIPHERTEXT_WIDTH'd9930709;
cipher_text[40] = `CIPHERTEXT_WIDTH'd9663207;
cipher_text[41] = `CIPHERTEXT_WIDTH'd12214005;
cipher_text[42] = `CIPHERTEXT_WIDTH'd6522228;
cipher_text[43] = `CIPHERTEXT_WIDTH'd1671125;
cipher_text[44] = `CIPHERTEXT_WIDTH'd3219493;
cipher_text[45] = `CIPHERTEXT_WIDTH'd2457812;
cipher_text[46] = `CIPHERTEXT_WIDTH'd10041809;
cipher_text[47] = `CIPHERTEXT_WIDTH'd1768975;
cipher_text[48] = `CIPHERTEXT_WIDTH'd12667909;
cipher_text[49] = `CIPHERTEXT_WIDTH'd7572873;
cipher_text[50] = `CIPHERTEXT_WIDTH'd3292911;
cipher_text[51] = `CIPHERTEXT_WIDTH'd11167755;
cipher_text[52] = `CIPHERTEXT_WIDTH'd1550567;
cipher_text[53] = `CIPHERTEXT_WIDTH'd7870366;
cipher_text[54] = `CIPHERTEXT_WIDTH'd5600744;
cipher_text[55] = `CIPHERTEXT_WIDTH'd2117351;
cipher_text[56] = `CIPHERTEXT_WIDTH'd229554;
cipher_text[57] = `CIPHERTEXT_WIDTH'd7436074;
cipher_text[58] = `CIPHERTEXT_WIDTH'd373030;
cipher_text[59] = `CIPHERTEXT_WIDTH'd1551185;
cipher_text[60] = `CIPHERTEXT_WIDTH'd5436356;
cipher_text[61] = `CIPHERTEXT_WIDTH'd9888525;
cipher_text[62] = `CIPHERTEXT_WIDTH'd8157063;
cipher_text[63] = `CIPHERTEXT_WIDTH'd1020403;
cipher_text[64] = `CIPHERTEXT_WIDTH'd12207997;
cipher_text[65] = `CIPHERTEXT_WIDTH'd1633388;
cipher_text[66] = `CIPHERTEXT_WIDTH'd12626307;
cipher_text[67] = `CIPHERTEXT_WIDTH'd15737951;
cipher_text[68] = `CIPHERTEXT_WIDTH'd2136404;
cipher_text[69] = `CIPHERTEXT_WIDTH'd2277438;
cipher_text[70] = `CIPHERTEXT_WIDTH'd3072190;
cipher_text[71] = `CIPHERTEXT_WIDTH'd12551248;
cipher_text[72] = `CIPHERTEXT_WIDTH'd1846568;
cipher_text[73] = `CIPHERTEXT_WIDTH'd3770541;
cipher_text[74] = `CIPHERTEXT_WIDTH'd13192398;
cipher_text[75] = `CIPHERTEXT_WIDTH'd16193154;
cipher_text[76] = `CIPHERTEXT_WIDTH'd5616110;
cipher_text[77] = `CIPHERTEXT_WIDTH'd14099700;
cipher_text[78] = `CIPHERTEXT_WIDTH'd10529371;
cipher_text[79] = `CIPHERTEXT_WIDTH'd1613472;
cipher_text[80] = `CIPHERTEXT_WIDTH'd14106904;
cipher_text[81] = `CIPHERTEXT_WIDTH'd16116559;
cipher_text[82] = `CIPHERTEXT_WIDTH'd9038126;
cipher_text[83] = `CIPHERTEXT_WIDTH'd7023256;
cipher_text[84] = `CIPHERTEXT_WIDTH'd15652169;
cipher_text[85] = `CIPHERTEXT_WIDTH'd6739754;
cipher_text[86] = `CIPHERTEXT_WIDTH'd3009580;
cipher_text[87] = `CIPHERTEXT_WIDTH'd10392477;
cipher_text[88] = `CIPHERTEXT_WIDTH'd15064007;
cipher_text[89] = `CIPHERTEXT_WIDTH'd16243582;
cipher_text[90] = `CIPHERTEXT_WIDTH'd903507;
cipher_text[91] = `CIPHERTEXT_WIDTH'd5430041;
cipher_text[92] = `CIPHERTEXT_WIDTH'd12304368;
cipher_text[93] = `CIPHERTEXT_WIDTH'd8087275;
cipher_text[94] = `CIPHERTEXT_WIDTH'd9476563;
cipher_text[95] = `CIPHERTEXT_WIDTH'd3853370;
cipher_text[96] = `CIPHERTEXT_WIDTH'd14818868;
cipher_text[97] = `CIPHERTEXT_WIDTH'd10402598;
cipher_text[98] = `CIPHERTEXT_WIDTH'd6709706;
cipher_text[99] = `CIPHERTEXT_WIDTH'd4377074;
cipher_text[100] = `CIPHERTEXT_WIDTH'd10760206;
cipher_text[101] = `CIPHERTEXT_WIDTH'd2060086;
cipher_text[102] = `CIPHERTEXT_WIDTH'd11959282;
cipher_text[103] = `CIPHERTEXT_WIDTH'd13473305;
cipher_text[104] = `CIPHERTEXT_WIDTH'd4196759;
cipher_text[105] = `CIPHERTEXT_WIDTH'd7541139;
cipher_text[106] = `CIPHERTEXT_WIDTH'd6331316;
cipher_text[107] = `CIPHERTEXT_WIDTH'd11552325;
cipher_text[108] = `CIPHERTEXT_WIDTH'd15787500;
cipher_text[109] = `CIPHERTEXT_WIDTH'd11117840;
cipher_text[110] = `CIPHERTEXT_WIDTH'd11817391;
cipher_text[111] = `CIPHERTEXT_WIDTH'd3619545;
cipher_text[112] = `CIPHERTEXT_WIDTH'd4974894;
cipher_text[113] = `CIPHERTEXT_WIDTH'd9912651;
cipher_text[114] = `CIPHERTEXT_WIDTH'd16491851;
cipher_text[115] = `CIPHERTEXT_WIDTH'd15798715;
cipher_text[116] = `CIPHERTEXT_WIDTH'd6486937;
cipher_text[117] = `CIPHERTEXT_WIDTH'd6342758;
cipher_text[118] = `CIPHERTEXT_WIDTH'd13044667;
cipher_text[119] = `CIPHERTEXT_WIDTH'd6716693;
cipher_text[120] = `CIPHERTEXT_WIDTH'd9465012;
cipher_text[121] = `CIPHERTEXT_WIDTH'd8547744;
cipher_text[122] = `CIPHERTEXT_WIDTH'd15574173;
cipher_text[123] = `CIPHERTEXT_WIDTH'd9595969;
cipher_text[124] = `CIPHERTEXT_WIDTH'd10605705;
cipher_text[125] = `CIPHERTEXT_WIDTH'd8537730;
cipher_text[126] = `CIPHERTEXT_WIDTH'd15081762;
cipher_text[127] = `CIPHERTEXT_WIDTH'd15000695;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 8;
cipher_text[0] = `CIPHERTEXT_WIDTH'd1165476;
cipher_text[1] = `CIPHERTEXT_WIDTH'd2716295;
cipher_text[2] = `CIPHERTEXT_WIDTH'd4258534;
cipher_text[3] = `CIPHERTEXT_WIDTH'd13008414;
cipher_text[4] = `CIPHERTEXT_WIDTH'd15238817;
cipher_text[5] = `CIPHERTEXT_WIDTH'd10228726;
cipher_text[6] = `CIPHERTEXT_WIDTH'd3920633;
cipher_text[7] = `CIPHERTEXT_WIDTH'd7294649;
cipher_text[8] = `CIPHERTEXT_WIDTH'd11823134;
cipher_text[9] = `CIPHERTEXT_WIDTH'd2966933;
cipher_text[10] = `CIPHERTEXT_WIDTH'd6304202;
cipher_text[11] = `CIPHERTEXT_WIDTH'd6559492;
cipher_text[12] = `CIPHERTEXT_WIDTH'd7332624;
cipher_text[13] = `CIPHERTEXT_WIDTH'd6307408;
cipher_text[14] = `CIPHERTEXT_WIDTH'd16381980;
cipher_text[15] = `CIPHERTEXT_WIDTH'd12819810;
cipher_text[16] = `CIPHERTEXT_WIDTH'd9968949;
cipher_text[17] = `CIPHERTEXT_WIDTH'd16182105;
cipher_text[18] = `CIPHERTEXT_WIDTH'd15918083;
cipher_text[19] = `CIPHERTEXT_WIDTH'd4315182;
cipher_text[20] = `CIPHERTEXT_WIDTH'd8562570;
cipher_text[21] = `CIPHERTEXT_WIDTH'd11887183;
cipher_text[22] = `CIPHERTEXT_WIDTH'd6897690;
cipher_text[23] = `CIPHERTEXT_WIDTH'd13226932;
cipher_text[24] = `CIPHERTEXT_WIDTH'd14587880;
cipher_text[25] = `CIPHERTEXT_WIDTH'd9014547;
cipher_text[26] = `CIPHERTEXT_WIDTH'd10233707;
cipher_text[27] = `CIPHERTEXT_WIDTH'd16699174;
cipher_text[28] = `CIPHERTEXT_WIDTH'd10596698;
cipher_text[29] = `CIPHERTEXT_WIDTH'd5053630;
cipher_text[30] = `CIPHERTEXT_WIDTH'd15046131;
cipher_text[31] = `CIPHERTEXT_WIDTH'd11950795;
cipher_text[32] = `CIPHERTEXT_WIDTH'd15741282;
cipher_text[33] = `CIPHERTEXT_WIDTH'd12785059;
cipher_text[34] = `CIPHERTEXT_WIDTH'd14900094;
cipher_text[35] = `CIPHERTEXT_WIDTH'd1143743;
cipher_text[36] = `CIPHERTEXT_WIDTH'd14731348;
cipher_text[37] = `CIPHERTEXT_WIDTH'd7339171;
cipher_text[38] = `CIPHERTEXT_WIDTH'd8403336;
cipher_text[39] = `CIPHERTEXT_WIDTH'd13966001;
cipher_text[40] = `CIPHERTEXT_WIDTH'd15015337;
cipher_text[41] = `CIPHERTEXT_WIDTH'd6022565;
cipher_text[42] = `CIPHERTEXT_WIDTH'd988453;
cipher_text[43] = `CIPHERTEXT_WIDTH'd9348731;
cipher_text[44] = `CIPHERTEXT_WIDTH'd8144435;
cipher_text[45] = `CIPHERTEXT_WIDTH'd1638099;
cipher_text[46] = `CIPHERTEXT_WIDTH'd13893557;
cipher_text[47] = `CIPHERTEXT_WIDTH'd4743418;
cipher_text[48] = `CIPHERTEXT_WIDTH'd2083858;
cipher_text[49] = `CIPHERTEXT_WIDTH'd9173782;
cipher_text[50] = `CIPHERTEXT_WIDTH'd993754;
cipher_text[51] = `CIPHERTEXT_WIDTH'd7758493;
cipher_text[52] = `CIPHERTEXT_WIDTH'd4832774;
cipher_text[53] = `CIPHERTEXT_WIDTH'd16272063;
cipher_text[54] = `CIPHERTEXT_WIDTH'd6057923;
cipher_text[55] = `CIPHERTEXT_WIDTH'd4433863;
cipher_text[56] = `CIPHERTEXT_WIDTH'd7954147;
cipher_text[57] = `CIPHERTEXT_WIDTH'd10230381;
cipher_text[58] = `CIPHERTEXT_WIDTH'd7350589;
cipher_text[59] = `CIPHERTEXT_WIDTH'd4628739;
cipher_text[60] = `CIPHERTEXT_WIDTH'd7974048;
cipher_text[61] = `CIPHERTEXT_WIDTH'd11844105;
cipher_text[62] = `CIPHERTEXT_WIDTH'd13163966;
cipher_text[63] = `CIPHERTEXT_WIDTH'd16355738;
cipher_text[64] = `CIPHERTEXT_WIDTH'd9021289;
cipher_text[65] = `CIPHERTEXT_WIDTH'd213115;
cipher_text[66] = `CIPHERTEXT_WIDTH'd4396415;
cipher_text[67] = `CIPHERTEXT_WIDTH'd12069134;
cipher_text[68] = `CIPHERTEXT_WIDTH'd515169;
cipher_text[69] = `CIPHERTEXT_WIDTH'd9368972;
cipher_text[70] = `CIPHERTEXT_WIDTH'd16133709;
cipher_text[71] = `CIPHERTEXT_WIDTH'd6774580;
cipher_text[72] = `CIPHERTEXT_WIDTH'd2360136;
cipher_text[73] = `CIPHERTEXT_WIDTH'd578096;
cipher_text[74] = `CIPHERTEXT_WIDTH'd3888258;
cipher_text[75] = `CIPHERTEXT_WIDTH'd13158632;
cipher_text[76] = `CIPHERTEXT_WIDTH'd5020292;
cipher_text[77] = `CIPHERTEXT_WIDTH'd926855;
cipher_text[78] = `CIPHERTEXT_WIDTH'd6466442;
cipher_text[79] = `CIPHERTEXT_WIDTH'd12131259;
cipher_text[80] = `CIPHERTEXT_WIDTH'd5617266;
cipher_text[81] = `CIPHERTEXT_WIDTH'd15281033;
cipher_text[82] = `CIPHERTEXT_WIDTH'd7937270;
cipher_text[83] = `CIPHERTEXT_WIDTH'd10934914;
cipher_text[84] = `CIPHERTEXT_WIDTH'd11591561;
cipher_text[85] = `CIPHERTEXT_WIDTH'd6199457;
cipher_text[86] = `CIPHERTEXT_WIDTH'd7883951;
cipher_text[87] = `CIPHERTEXT_WIDTH'd12758959;
cipher_text[88] = `CIPHERTEXT_WIDTH'd9314918;
cipher_text[89] = `CIPHERTEXT_WIDTH'd4943762;
cipher_text[90] = `CIPHERTEXT_WIDTH'd13700765;
cipher_text[91] = `CIPHERTEXT_WIDTH'd10590490;
cipher_text[92] = `CIPHERTEXT_WIDTH'd5033998;
cipher_text[93] = `CIPHERTEXT_WIDTH'd4850186;
cipher_text[94] = `CIPHERTEXT_WIDTH'd9878707;
cipher_text[95] = `CIPHERTEXT_WIDTH'd7949613;
cipher_text[96] = `CIPHERTEXT_WIDTH'd15209063;
cipher_text[97] = `CIPHERTEXT_WIDTH'd9556844;
cipher_text[98] = `CIPHERTEXT_WIDTH'd5782650;
cipher_text[99] = `CIPHERTEXT_WIDTH'd4446233;
cipher_text[100] = `CIPHERTEXT_WIDTH'd10776310;
cipher_text[101] = `CIPHERTEXT_WIDTH'd8608542;
cipher_text[102] = `CIPHERTEXT_WIDTH'd5116130;
cipher_text[103] = `CIPHERTEXT_WIDTH'd4405870;
cipher_text[104] = `CIPHERTEXT_WIDTH'd8211583;
cipher_text[105] = `CIPHERTEXT_WIDTH'd13473710;
cipher_text[106] = `CIPHERTEXT_WIDTH'd9767296;
cipher_text[107] = `CIPHERTEXT_WIDTH'd6403937;
cipher_text[108] = `CIPHERTEXT_WIDTH'd1994565;
cipher_text[109] = `CIPHERTEXT_WIDTH'd1978592;
cipher_text[110] = `CIPHERTEXT_WIDTH'd13015090;
cipher_text[111] = `CIPHERTEXT_WIDTH'd6243962;
cipher_text[112] = `CIPHERTEXT_WIDTH'd11993221;
cipher_text[113] = `CIPHERTEXT_WIDTH'd894486;
cipher_text[114] = `CIPHERTEXT_WIDTH'd11017432;
cipher_text[115] = `CIPHERTEXT_WIDTH'd11654238;
cipher_text[116] = `CIPHERTEXT_WIDTH'd13362616;
cipher_text[117] = `CIPHERTEXT_WIDTH'd6041685;
cipher_text[118] = `CIPHERTEXT_WIDTH'd11369755;
cipher_text[119] = `CIPHERTEXT_WIDTH'd14962968;
cipher_text[120] = `CIPHERTEXT_WIDTH'd3153505;
cipher_text[121] = `CIPHERTEXT_WIDTH'd12558994;
cipher_text[122] = `CIPHERTEXT_WIDTH'd16724330;
cipher_text[123] = `CIPHERTEXT_WIDTH'd5641823;
cipher_text[124] = `CIPHERTEXT_WIDTH'd5556793;
cipher_text[125] = `CIPHERTEXT_WIDTH'd388774;
cipher_text[126] = `CIPHERTEXT_WIDTH'd2981719;
cipher_text[127] = `CIPHERTEXT_WIDTH'd7665932;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 9;
cipher_text[0] = `CIPHERTEXT_WIDTH'd13452497;
cipher_text[1] = `CIPHERTEXT_WIDTH'd4160083;
cipher_text[2] = `CIPHERTEXT_WIDTH'd16340316;
cipher_text[3] = `CIPHERTEXT_WIDTH'd15312652;
cipher_text[4] = `CIPHERTEXT_WIDTH'd14274758;
cipher_text[5] = `CIPHERTEXT_WIDTH'd141232;
cipher_text[6] = `CIPHERTEXT_WIDTH'd3219427;
cipher_text[7] = `CIPHERTEXT_WIDTH'd7787671;
cipher_text[8] = `CIPHERTEXT_WIDTH'd11851388;
cipher_text[9] = `CIPHERTEXT_WIDTH'd12986125;
cipher_text[10] = `CIPHERTEXT_WIDTH'd358937;
cipher_text[11] = `CIPHERTEXT_WIDTH'd11226328;
cipher_text[12] = `CIPHERTEXT_WIDTH'd10563288;
cipher_text[13] = `CIPHERTEXT_WIDTH'd1824122;
cipher_text[14] = `CIPHERTEXT_WIDTH'd7007791;
cipher_text[15] = `CIPHERTEXT_WIDTH'd12227666;
cipher_text[16] = `CIPHERTEXT_WIDTH'd8092845;
cipher_text[17] = `CIPHERTEXT_WIDTH'd15603754;
cipher_text[18] = `CIPHERTEXT_WIDTH'd4775847;
cipher_text[19] = `CIPHERTEXT_WIDTH'd9009226;
cipher_text[20] = `CIPHERTEXT_WIDTH'd5972583;
cipher_text[21] = `CIPHERTEXT_WIDTH'd5779587;
cipher_text[22] = `CIPHERTEXT_WIDTH'd11355950;
cipher_text[23] = `CIPHERTEXT_WIDTH'd9914243;
cipher_text[24] = `CIPHERTEXT_WIDTH'd3211578;
cipher_text[25] = `CIPHERTEXT_WIDTH'd16383042;
cipher_text[26] = `CIPHERTEXT_WIDTH'd6615167;
cipher_text[27] = `CIPHERTEXT_WIDTH'd3258955;
cipher_text[28] = `CIPHERTEXT_WIDTH'd13994828;
cipher_text[29] = `CIPHERTEXT_WIDTH'd4090900;
cipher_text[30] = `CIPHERTEXT_WIDTH'd4565875;
cipher_text[31] = `CIPHERTEXT_WIDTH'd15624968;
cipher_text[32] = `CIPHERTEXT_WIDTH'd14048160;
cipher_text[33] = `CIPHERTEXT_WIDTH'd4984040;
cipher_text[34] = `CIPHERTEXT_WIDTH'd7639009;
cipher_text[35] = `CIPHERTEXT_WIDTH'd5860652;
cipher_text[36] = `CIPHERTEXT_WIDTH'd2050987;
cipher_text[37] = `CIPHERTEXT_WIDTH'd12006654;
cipher_text[38] = `CIPHERTEXT_WIDTH'd3185569;
cipher_text[39] = `CIPHERTEXT_WIDTH'd5073846;
cipher_text[40] = `CIPHERTEXT_WIDTH'd13688855;
cipher_text[41] = `CIPHERTEXT_WIDTH'd12758285;
cipher_text[42] = `CIPHERTEXT_WIDTH'd12088671;
cipher_text[43] = `CIPHERTEXT_WIDTH'd7893556;
cipher_text[44] = `CIPHERTEXT_WIDTH'd11411458;
cipher_text[45] = `CIPHERTEXT_WIDTH'd16711316;
cipher_text[46] = `CIPHERTEXT_WIDTH'd9714881;
cipher_text[47] = `CIPHERTEXT_WIDTH'd3178071;
cipher_text[48] = `CIPHERTEXT_WIDTH'd10903907;
cipher_text[49] = `CIPHERTEXT_WIDTH'd8473077;
cipher_text[50] = `CIPHERTEXT_WIDTH'd5405214;
cipher_text[51] = `CIPHERTEXT_WIDTH'd11969406;
cipher_text[52] = `CIPHERTEXT_WIDTH'd10648220;
cipher_text[53] = `CIPHERTEXT_WIDTH'd5357877;
cipher_text[54] = `CIPHERTEXT_WIDTH'd12186604;
cipher_text[55] = `CIPHERTEXT_WIDTH'd16565618;
cipher_text[56] = `CIPHERTEXT_WIDTH'd15215429;
cipher_text[57] = `CIPHERTEXT_WIDTH'd4202644;
cipher_text[58] = `CIPHERTEXT_WIDTH'd6947090;
cipher_text[59] = `CIPHERTEXT_WIDTH'd12929073;
cipher_text[60] = `CIPHERTEXT_WIDTH'd10143836;
cipher_text[61] = `CIPHERTEXT_WIDTH'd14668623;
cipher_text[62] = `CIPHERTEXT_WIDTH'd7129951;
cipher_text[63] = `CIPHERTEXT_WIDTH'd5816242;
cipher_text[64] = `CIPHERTEXT_WIDTH'd5325028;
cipher_text[65] = `CIPHERTEXT_WIDTH'd7930046;
cipher_text[66] = `CIPHERTEXT_WIDTH'd10017781;
cipher_text[67] = `CIPHERTEXT_WIDTH'd1098925;
cipher_text[68] = `CIPHERTEXT_WIDTH'd6592495;
cipher_text[69] = `CIPHERTEXT_WIDTH'd10365854;
cipher_text[70] = `CIPHERTEXT_WIDTH'd11047690;
cipher_text[71] = `CIPHERTEXT_WIDTH'd16452249;
cipher_text[72] = `CIPHERTEXT_WIDTH'd9890651;
cipher_text[73] = `CIPHERTEXT_WIDTH'd4898346;
cipher_text[74] = `CIPHERTEXT_WIDTH'd425939;
cipher_text[75] = `CIPHERTEXT_WIDTH'd10351014;
cipher_text[76] = `CIPHERTEXT_WIDTH'd11548173;
cipher_text[77] = `CIPHERTEXT_WIDTH'd12958879;
cipher_text[78] = `CIPHERTEXT_WIDTH'd9144000;
cipher_text[79] = `CIPHERTEXT_WIDTH'd12024583;
cipher_text[80] = `CIPHERTEXT_WIDTH'd15319530;
cipher_text[81] = `CIPHERTEXT_WIDTH'd16225857;
cipher_text[82] = `CIPHERTEXT_WIDTH'd5137654;
cipher_text[83] = `CIPHERTEXT_WIDTH'd1073228;
cipher_text[84] = `CIPHERTEXT_WIDTH'd14988497;
cipher_text[85] = `CIPHERTEXT_WIDTH'd430349;
cipher_text[86] = `CIPHERTEXT_WIDTH'd10043398;
cipher_text[87] = `CIPHERTEXT_WIDTH'd7827992;
cipher_text[88] = `CIPHERTEXT_WIDTH'd15717419;
cipher_text[89] = `CIPHERTEXT_WIDTH'd1086874;
cipher_text[90] = `CIPHERTEXT_WIDTH'd8788979;
cipher_text[91] = `CIPHERTEXT_WIDTH'd7312304;
cipher_text[92] = `CIPHERTEXT_WIDTH'd12517371;
cipher_text[93] = `CIPHERTEXT_WIDTH'd7887307;
cipher_text[94] = `CIPHERTEXT_WIDTH'd11354557;
cipher_text[95] = `CIPHERTEXT_WIDTH'd13288955;
cipher_text[96] = `CIPHERTEXT_WIDTH'd10216736;
cipher_text[97] = `CIPHERTEXT_WIDTH'd8429506;
cipher_text[98] = `CIPHERTEXT_WIDTH'd10516058;
cipher_text[99] = `CIPHERTEXT_WIDTH'd981657;
cipher_text[100] = `CIPHERTEXT_WIDTH'd4988044;
cipher_text[101] = `CIPHERTEXT_WIDTH'd14086727;
cipher_text[102] = `CIPHERTEXT_WIDTH'd6634472;
cipher_text[103] = `CIPHERTEXT_WIDTH'd10614009;
cipher_text[104] = `CIPHERTEXT_WIDTH'd9399986;
cipher_text[105] = `CIPHERTEXT_WIDTH'd368303;
cipher_text[106] = `CIPHERTEXT_WIDTH'd2642875;
cipher_text[107] = `CIPHERTEXT_WIDTH'd7569708;
cipher_text[108] = `CIPHERTEXT_WIDTH'd10057501;
cipher_text[109] = `CIPHERTEXT_WIDTH'd9883714;
cipher_text[110] = `CIPHERTEXT_WIDTH'd178890;
cipher_text[111] = `CIPHERTEXT_WIDTH'd746617;
cipher_text[112] = `CIPHERTEXT_WIDTH'd15934229;
cipher_text[113] = `CIPHERTEXT_WIDTH'd11027872;
cipher_text[114] = `CIPHERTEXT_WIDTH'd10116339;
cipher_text[115] = `CIPHERTEXT_WIDTH'd15936775;
cipher_text[116] = `CIPHERTEXT_WIDTH'd1941374;
cipher_text[117] = `CIPHERTEXT_WIDTH'd2009370;
cipher_text[118] = `CIPHERTEXT_WIDTH'd7579875;
cipher_text[119] = `CIPHERTEXT_WIDTH'd1009151;
cipher_text[120] = `CIPHERTEXT_WIDTH'd3639792;
cipher_text[121] = `CIPHERTEXT_WIDTH'd6376162;
cipher_text[122] = `CIPHERTEXT_WIDTH'd12984659;
cipher_text[123] = `CIPHERTEXT_WIDTH'd7349773;
cipher_text[124] = `CIPHERTEXT_WIDTH'd9588214;
cipher_text[125] = `CIPHERTEXT_WIDTH'd10550410;
cipher_text[126] = `CIPHERTEXT_WIDTH'd8291191;
cipher_text[127] = `CIPHERTEXT_WIDTH'd850037;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 10;
cipher_text[0] = `CIPHERTEXT_WIDTH'd15123380;
cipher_text[1] = `CIPHERTEXT_WIDTH'd574355;
cipher_text[2] = `CIPHERTEXT_WIDTH'd14339286;
cipher_text[3] = `CIPHERTEXT_WIDTH'd4799826;
cipher_text[4] = `CIPHERTEXT_WIDTH'd11208796;
cipher_text[5] = `CIPHERTEXT_WIDTH'd10882925;
cipher_text[6] = `CIPHERTEXT_WIDTH'd9108497;
cipher_text[7] = `CIPHERTEXT_WIDTH'd16302507;
cipher_text[8] = `CIPHERTEXT_WIDTH'd4444079;
cipher_text[9] = `CIPHERTEXT_WIDTH'd4120009;
cipher_text[10] = `CIPHERTEXT_WIDTH'd14579135;
cipher_text[11] = `CIPHERTEXT_WIDTH'd2886436;
cipher_text[12] = `CIPHERTEXT_WIDTH'd5409789;
cipher_text[13] = `CIPHERTEXT_WIDTH'd11713773;
cipher_text[14] = `CIPHERTEXT_WIDTH'd7634454;
cipher_text[15] = `CIPHERTEXT_WIDTH'd4650784;
cipher_text[16] = `CIPHERTEXT_WIDTH'd239378;
cipher_text[17] = `CIPHERTEXT_WIDTH'd7403993;
cipher_text[18] = `CIPHERTEXT_WIDTH'd16033908;
cipher_text[19] = `CIPHERTEXT_WIDTH'd6363837;
cipher_text[20] = `CIPHERTEXT_WIDTH'd3751536;
cipher_text[21] = `CIPHERTEXT_WIDTH'd10824003;
cipher_text[22] = `CIPHERTEXT_WIDTH'd14084316;
cipher_text[23] = `CIPHERTEXT_WIDTH'd12666336;
cipher_text[24] = `CIPHERTEXT_WIDTH'd11335843;
cipher_text[25] = `CIPHERTEXT_WIDTH'd7546607;
cipher_text[26] = `CIPHERTEXT_WIDTH'd12033027;
cipher_text[27] = `CIPHERTEXT_WIDTH'd6305295;
cipher_text[28] = `CIPHERTEXT_WIDTH'd9127247;
cipher_text[29] = `CIPHERTEXT_WIDTH'd5848741;
cipher_text[30] = `CIPHERTEXT_WIDTH'd4864443;
cipher_text[31] = `CIPHERTEXT_WIDTH'd16678716;
cipher_text[32] = `CIPHERTEXT_WIDTH'd4780907;
cipher_text[33] = `CIPHERTEXT_WIDTH'd7707340;
cipher_text[34] = `CIPHERTEXT_WIDTH'd10511537;
cipher_text[35] = `CIPHERTEXT_WIDTH'd10661329;
cipher_text[36] = `CIPHERTEXT_WIDTH'd15149069;
cipher_text[37] = `CIPHERTEXT_WIDTH'd5182568;
cipher_text[38] = `CIPHERTEXT_WIDTH'd5352699;
cipher_text[39] = `CIPHERTEXT_WIDTH'd394603;
cipher_text[40] = `CIPHERTEXT_WIDTH'd8618603;
cipher_text[41] = `CIPHERTEXT_WIDTH'd11024180;
cipher_text[42] = `CIPHERTEXT_WIDTH'd12376177;
cipher_text[43] = `CIPHERTEXT_WIDTH'd7439684;
cipher_text[44] = `CIPHERTEXT_WIDTH'd13945546;
cipher_text[45] = `CIPHERTEXT_WIDTH'd15833931;
cipher_text[46] = `CIPHERTEXT_WIDTH'd1626727;
cipher_text[47] = `CIPHERTEXT_WIDTH'd15057113;
cipher_text[48] = `CIPHERTEXT_WIDTH'd9535928;
cipher_text[49] = `CIPHERTEXT_WIDTH'd5286336;
cipher_text[50] = `CIPHERTEXT_WIDTH'd12711921;
cipher_text[51] = `CIPHERTEXT_WIDTH'd314392;
cipher_text[52] = `CIPHERTEXT_WIDTH'd2448596;
cipher_text[53] = `CIPHERTEXT_WIDTH'd4164470;
cipher_text[54] = `CIPHERTEXT_WIDTH'd6509954;
cipher_text[55] = `CIPHERTEXT_WIDTH'd11504794;
cipher_text[56] = `CIPHERTEXT_WIDTH'd15768187;
cipher_text[57] = `CIPHERTEXT_WIDTH'd3373634;
cipher_text[58] = `CIPHERTEXT_WIDTH'd645016;
cipher_text[59] = `CIPHERTEXT_WIDTH'd4106276;
cipher_text[60] = `CIPHERTEXT_WIDTH'd16390882;
cipher_text[61] = `CIPHERTEXT_WIDTH'd9195614;
cipher_text[62] = `CIPHERTEXT_WIDTH'd12485823;
cipher_text[63] = `CIPHERTEXT_WIDTH'd9893044;
cipher_text[64] = `CIPHERTEXT_WIDTH'd14171913;
cipher_text[65] = `CIPHERTEXT_WIDTH'd4071517;
cipher_text[66] = `CIPHERTEXT_WIDTH'd12955978;
cipher_text[67] = `CIPHERTEXT_WIDTH'd12240974;
cipher_text[68] = `CIPHERTEXT_WIDTH'd15534924;
cipher_text[69] = `CIPHERTEXT_WIDTH'd776272;
cipher_text[70] = `CIPHERTEXT_WIDTH'd11538717;
cipher_text[71] = `CIPHERTEXT_WIDTH'd4848024;
cipher_text[72] = `CIPHERTEXT_WIDTH'd12945198;
cipher_text[73] = `CIPHERTEXT_WIDTH'd5535697;
cipher_text[74] = `CIPHERTEXT_WIDTH'd16488900;
cipher_text[75] = `CIPHERTEXT_WIDTH'd13678535;
cipher_text[76] = `CIPHERTEXT_WIDTH'd7552003;
cipher_text[77] = `CIPHERTEXT_WIDTH'd10689427;
cipher_text[78] = `CIPHERTEXT_WIDTH'd11871501;
cipher_text[79] = `CIPHERTEXT_WIDTH'd6286901;
cipher_text[80] = `CIPHERTEXT_WIDTH'd9233692;
cipher_text[81] = `CIPHERTEXT_WIDTH'd10540923;
cipher_text[82] = `CIPHERTEXT_WIDTH'd8584715;
cipher_text[83] = `CIPHERTEXT_WIDTH'd2545343;
cipher_text[84] = `CIPHERTEXT_WIDTH'd9350512;
cipher_text[85] = `CIPHERTEXT_WIDTH'd15958833;
cipher_text[86] = `CIPHERTEXT_WIDTH'd14726765;
cipher_text[87] = `CIPHERTEXT_WIDTH'd6305534;
cipher_text[88] = `CIPHERTEXT_WIDTH'd10116713;
cipher_text[89] = `CIPHERTEXT_WIDTH'd8895224;
cipher_text[90] = `CIPHERTEXT_WIDTH'd12817555;
cipher_text[91] = `CIPHERTEXT_WIDTH'd8923429;
cipher_text[92] = `CIPHERTEXT_WIDTH'd1319367;
cipher_text[93] = `CIPHERTEXT_WIDTH'd11830742;
cipher_text[94] = `CIPHERTEXT_WIDTH'd14394777;
cipher_text[95] = `CIPHERTEXT_WIDTH'd6706804;
cipher_text[96] = `CIPHERTEXT_WIDTH'd1503235;
cipher_text[97] = `CIPHERTEXT_WIDTH'd568007;
cipher_text[98] = `CIPHERTEXT_WIDTH'd13017521;
cipher_text[99] = `CIPHERTEXT_WIDTH'd14903384;
cipher_text[100] = `CIPHERTEXT_WIDTH'd9685512;
cipher_text[101] = `CIPHERTEXT_WIDTH'd15074694;
cipher_text[102] = `CIPHERTEXT_WIDTH'd9779746;
cipher_text[103] = `CIPHERTEXT_WIDTH'd3211113;
cipher_text[104] = `CIPHERTEXT_WIDTH'd10381289;
cipher_text[105] = `CIPHERTEXT_WIDTH'd2326290;
cipher_text[106] = `CIPHERTEXT_WIDTH'd10332488;
cipher_text[107] = `CIPHERTEXT_WIDTH'd6097037;
cipher_text[108] = `CIPHERTEXT_WIDTH'd14166846;
cipher_text[109] = `CIPHERTEXT_WIDTH'd206247;
cipher_text[110] = `CIPHERTEXT_WIDTH'd15077521;
cipher_text[111] = `CIPHERTEXT_WIDTH'd2120073;
cipher_text[112] = `CIPHERTEXT_WIDTH'd6839895;
cipher_text[113] = `CIPHERTEXT_WIDTH'd13748972;
cipher_text[114] = `CIPHERTEXT_WIDTH'd7250688;
cipher_text[115] = `CIPHERTEXT_WIDTH'd16281603;
cipher_text[116] = `CIPHERTEXT_WIDTH'd13172148;
cipher_text[117] = `CIPHERTEXT_WIDTH'd14505736;
cipher_text[118] = `CIPHERTEXT_WIDTH'd4563655;
cipher_text[119] = `CIPHERTEXT_WIDTH'd11809837;
cipher_text[120] = `CIPHERTEXT_WIDTH'd3651064;
cipher_text[121] = `CIPHERTEXT_WIDTH'd11475780;
cipher_text[122] = `CIPHERTEXT_WIDTH'd7945919;
cipher_text[123] = `CIPHERTEXT_WIDTH'd15919779;
cipher_text[124] = `CIPHERTEXT_WIDTH'd623186;
cipher_text[125] = `CIPHERTEXT_WIDTH'd9083756;
cipher_text[126] = `CIPHERTEXT_WIDTH'd1884494;
cipher_text[127] = `CIPHERTEXT_WIDTH'd4984032;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 11;
cipher_text[0] = `CIPHERTEXT_WIDTH'd6316762;
cipher_text[1] = `CIPHERTEXT_WIDTH'd10914157;
cipher_text[2] = `CIPHERTEXT_WIDTH'd1493722;
cipher_text[3] = `CIPHERTEXT_WIDTH'd10487196;
cipher_text[4] = `CIPHERTEXT_WIDTH'd10706190;
cipher_text[5] = `CIPHERTEXT_WIDTH'd1154066;
cipher_text[6] = `CIPHERTEXT_WIDTH'd2289847;
cipher_text[7] = `CIPHERTEXT_WIDTH'd12230545;
cipher_text[8] = `CIPHERTEXT_WIDTH'd5811439;
cipher_text[9] = `CIPHERTEXT_WIDTH'd15476593;
cipher_text[10] = `CIPHERTEXT_WIDTH'd5914334;
cipher_text[11] = `CIPHERTEXT_WIDTH'd1012843;
cipher_text[12] = `CIPHERTEXT_WIDTH'd14883107;
cipher_text[13] = `CIPHERTEXT_WIDTH'd4213510;
cipher_text[14] = `CIPHERTEXT_WIDTH'd3172115;
cipher_text[15] = `CIPHERTEXT_WIDTH'd11166851;
cipher_text[16] = `CIPHERTEXT_WIDTH'd4969022;
cipher_text[17] = `CIPHERTEXT_WIDTH'd4249282;
cipher_text[18] = `CIPHERTEXT_WIDTH'd3483855;
cipher_text[19] = `CIPHERTEXT_WIDTH'd2952064;
cipher_text[20] = `CIPHERTEXT_WIDTH'd5580229;
cipher_text[21] = `CIPHERTEXT_WIDTH'd9810577;
cipher_text[22] = `CIPHERTEXT_WIDTH'd5482271;
cipher_text[23] = `CIPHERTEXT_WIDTH'd4068660;
cipher_text[24] = `CIPHERTEXT_WIDTH'd3172729;
cipher_text[25] = `CIPHERTEXT_WIDTH'd10160606;
cipher_text[26] = `CIPHERTEXT_WIDTH'd14194050;
cipher_text[27] = `CIPHERTEXT_WIDTH'd9704143;
cipher_text[28] = `CIPHERTEXT_WIDTH'd13903015;
cipher_text[29] = `CIPHERTEXT_WIDTH'd811549;
cipher_text[30] = `CIPHERTEXT_WIDTH'd3635511;
cipher_text[31] = `CIPHERTEXT_WIDTH'd14651471;
cipher_text[32] = `CIPHERTEXT_WIDTH'd6936317;
cipher_text[33] = `CIPHERTEXT_WIDTH'd11623706;
cipher_text[34] = `CIPHERTEXT_WIDTH'd12265828;
cipher_text[35] = `CIPHERTEXT_WIDTH'd6844339;
cipher_text[36] = `CIPHERTEXT_WIDTH'd8258698;
cipher_text[37] = `CIPHERTEXT_WIDTH'd15396516;
cipher_text[38] = `CIPHERTEXT_WIDTH'd745845;
cipher_text[39] = `CIPHERTEXT_WIDTH'd14992123;
cipher_text[40] = `CIPHERTEXT_WIDTH'd12334639;
cipher_text[41] = `CIPHERTEXT_WIDTH'd9228308;
cipher_text[42] = `CIPHERTEXT_WIDTH'd4811901;
cipher_text[43] = `CIPHERTEXT_WIDTH'd3510608;
cipher_text[44] = `CIPHERTEXT_WIDTH'd15516830;
cipher_text[45] = `CIPHERTEXT_WIDTH'd170209;
cipher_text[46] = `CIPHERTEXT_WIDTH'd2592743;
cipher_text[47] = `CIPHERTEXT_WIDTH'd12839252;
cipher_text[48] = `CIPHERTEXT_WIDTH'd16673737;
cipher_text[49] = `CIPHERTEXT_WIDTH'd6180153;
cipher_text[50] = `CIPHERTEXT_WIDTH'd9981606;
cipher_text[51] = `CIPHERTEXT_WIDTH'd12322110;
cipher_text[52] = `CIPHERTEXT_WIDTH'd7605392;
cipher_text[53] = `CIPHERTEXT_WIDTH'd15963237;
cipher_text[54] = `CIPHERTEXT_WIDTH'd4994453;
cipher_text[55] = `CIPHERTEXT_WIDTH'd13353140;
cipher_text[56] = `CIPHERTEXT_WIDTH'd13126627;
cipher_text[57] = `CIPHERTEXT_WIDTH'd6718000;
cipher_text[58] = `CIPHERTEXT_WIDTH'd13672122;
cipher_text[59] = `CIPHERTEXT_WIDTH'd10825708;
cipher_text[60] = `CIPHERTEXT_WIDTH'd9936331;
cipher_text[61] = `CIPHERTEXT_WIDTH'd5424924;
cipher_text[62] = `CIPHERTEXT_WIDTH'd2393792;
cipher_text[63] = `CIPHERTEXT_WIDTH'd11086778;
cipher_text[64] = `CIPHERTEXT_WIDTH'd7625585;
cipher_text[65] = `CIPHERTEXT_WIDTH'd16260214;
cipher_text[66] = `CIPHERTEXT_WIDTH'd1197656;
cipher_text[67] = `CIPHERTEXT_WIDTH'd10766455;
cipher_text[68] = `CIPHERTEXT_WIDTH'd14085563;
cipher_text[69] = `CIPHERTEXT_WIDTH'd15664619;
cipher_text[70] = `CIPHERTEXT_WIDTH'd249275;
cipher_text[71] = `CIPHERTEXT_WIDTH'd6914953;
cipher_text[72] = `CIPHERTEXT_WIDTH'd7687314;
cipher_text[73] = `CIPHERTEXT_WIDTH'd2744873;
cipher_text[74] = `CIPHERTEXT_WIDTH'd13593911;
cipher_text[75] = `CIPHERTEXT_WIDTH'd457673;
cipher_text[76] = `CIPHERTEXT_WIDTH'd8431830;
cipher_text[77] = `CIPHERTEXT_WIDTH'd11627287;
cipher_text[78] = `CIPHERTEXT_WIDTH'd3428538;
cipher_text[79] = `CIPHERTEXT_WIDTH'd3264166;
cipher_text[80] = `CIPHERTEXT_WIDTH'd16491792;
cipher_text[81] = `CIPHERTEXT_WIDTH'd631149;
cipher_text[82] = `CIPHERTEXT_WIDTH'd6534177;
cipher_text[83] = `CIPHERTEXT_WIDTH'd14962673;
cipher_text[84] = `CIPHERTEXT_WIDTH'd11328235;
cipher_text[85] = `CIPHERTEXT_WIDTH'd3715185;
cipher_text[86] = `CIPHERTEXT_WIDTH'd4910979;
cipher_text[87] = `CIPHERTEXT_WIDTH'd14964215;
cipher_text[88] = `CIPHERTEXT_WIDTH'd5795375;
cipher_text[89] = `CIPHERTEXT_WIDTH'd7085620;
cipher_text[90] = `CIPHERTEXT_WIDTH'd8752760;
cipher_text[91] = `CIPHERTEXT_WIDTH'd12565105;
cipher_text[92] = `CIPHERTEXT_WIDTH'd5126294;
cipher_text[93] = `CIPHERTEXT_WIDTH'd10890152;
cipher_text[94] = `CIPHERTEXT_WIDTH'd6248675;
cipher_text[95] = `CIPHERTEXT_WIDTH'd7267947;
cipher_text[96] = `CIPHERTEXT_WIDTH'd15444438;
cipher_text[97] = `CIPHERTEXT_WIDTH'd6849467;
cipher_text[98] = `CIPHERTEXT_WIDTH'd6781735;
cipher_text[99] = `CIPHERTEXT_WIDTH'd9128238;
cipher_text[100] = `CIPHERTEXT_WIDTH'd759420;
cipher_text[101] = `CIPHERTEXT_WIDTH'd6634164;
cipher_text[102] = `CIPHERTEXT_WIDTH'd7751042;
cipher_text[103] = `CIPHERTEXT_WIDTH'd13445797;
cipher_text[104] = `CIPHERTEXT_WIDTH'd4351879;
cipher_text[105] = `CIPHERTEXT_WIDTH'd4589045;
cipher_text[106] = `CIPHERTEXT_WIDTH'd15309775;
cipher_text[107] = `CIPHERTEXT_WIDTH'd3434321;
cipher_text[108] = `CIPHERTEXT_WIDTH'd2362414;
cipher_text[109] = `CIPHERTEXT_WIDTH'd9506612;
cipher_text[110] = `CIPHERTEXT_WIDTH'd3503197;
cipher_text[111] = `CIPHERTEXT_WIDTH'd15063390;
cipher_text[112] = `CIPHERTEXT_WIDTH'd7809787;
cipher_text[113] = `CIPHERTEXT_WIDTH'd1234210;
cipher_text[114] = `CIPHERTEXT_WIDTH'd8726789;
cipher_text[115] = `CIPHERTEXT_WIDTH'd3365848;
cipher_text[116] = `CIPHERTEXT_WIDTH'd3198135;
cipher_text[117] = `CIPHERTEXT_WIDTH'd16364852;
cipher_text[118] = `CIPHERTEXT_WIDTH'd9504140;
cipher_text[119] = `CIPHERTEXT_WIDTH'd16662197;
cipher_text[120] = `CIPHERTEXT_WIDTH'd4262594;
cipher_text[121] = `CIPHERTEXT_WIDTH'd16600720;
cipher_text[122] = `CIPHERTEXT_WIDTH'd12279922;
cipher_text[123] = `CIPHERTEXT_WIDTH'd11897684;
cipher_text[124] = `CIPHERTEXT_WIDTH'd16101434;
cipher_text[125] = `CIPHERTEXT_WIDTH'd7814285;
cipher_text[126] = `CIPHERTEXT_WIDTH'd7554743;
cipher_text[127] = `CIPHERTEXT_WIDTH'd3163702;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 12;
cipher_text[0] = `CIPHERTEXT_WIDTH'd14040105;
cipher_text[1] = `CIPHERTEXT_WIDTH'd6458844;
cipher_text[2] = `CIPHERTEXT_WIDTH'd4574840;
cipher_text[3] = `CIPHERTEXT_WIDTH'd11906115;
cipher_text[4] = `CIPHERTEXT_WIDTH'd2185075;
cipher_text[5] = `CIPHERTEXT_WIDTH'd11931374;
cipher_text[6] = `CIPHERTEXT_WIDTH'd4618919;
cipher_text[7] = `CIPHERTEXT_WIDTH'd2282028;
cipher_text[8] = `CIPHERTEXT_WIDTH'd8050868;
cipher_text[9] = `CIPHERTEXT_WIDTH'd11900822;
cipher_text[10] = `CIPHERTEXT_WIDTH'd11902552;
cipher_text[11] = `CIPHERTEXT_WIDTH'd12368653;
cipher_text[12] = `CIPHERTEXT_WIDTH'd7488009;
cipher_text[13] = `CIPHERTEXT_WIDTH'd7433521;
cipher_text[14] = `CIPHERTEXT_WIDTH'd10340145;
cipher_text[15] = `CIPHERTEXT_WIDTH'd4393934;
cipher_text[16] = `CIPHERTEXT_WIDTH'd5900876;
cipher_text[17] = `CIPHERTEXT_WIDTH'd4246017;
cipher_text[18] = `CIPHERTEXT_WIDTH'd9520958;
cipher_text[19] = `CIPHERTEXT_WIDTH'd7366605;
cipher_text[20] = `CIPHERTEXT_WIDTH'd4074196;
cipher_text[21] = `CIPHERTEXT_WIDTH'd12036087;
cipher_text[22] = `CIPHERTEXT_WIDTH'd12148388;
cipher_text[23] = `CIPHERTEXT_WIDTH'd42449;
cipher_text[24] = `CIPHERTEXT_WIDTH'd2308664;
cipher_text[25] = `CIPHERTEXT_WIDTH'd3102696;
cipher_text[26] = `CIPHERTEXT_WIDTH'd16436405;
cipher_text[27] = `CIPHERTEXT_WIDTH'd1697460;
cipher_text[28] = `CIPHERTEXT_WIDTH'd4511213;
cipher_text[29] = `CIPHERTEXT_WIDTH'd11846295;
cipher_text[30] = `CIPHERTEXT_WIDTH'd15278897;
cipher_text[31] = `CIPHERTEXT_WIDTH'd8135802;
cipher_text[32] = `CIPHERTEXT_WIDTH'd6400781;
cipher_text[33] = `CIPHERTEXT_WIDTH'd13637131;
cipher_text[34] = `CIPHERTEXT_WIDTH'd13256711;
cipher_text[35] = `CIPHERTEXT_WIDTH'd13358237;
cipher_text[36] = `CIPHERTEXT_WIDTH'd7888600;
cipher_text[37] = `CIPHERTEXT_WIDTH'd11936520;
cipher_text[38] = `CIPHERTEXT_WIDTH'd12272748;
cipher_text[39] = `CIPHERTEXT_WIDTH'd13306211;
cipher_text[40] = `CIPHERTEXT_WIDTH'd4258652;
cipher_text[41] = `CIPHERTEXT_WIDTH'd11537281;
cipher_text[42] = `CIPHERTEXT_WIDTH'd8888429;
cipher_text[43] = `CIPHERTEXT_WIDTH'd7500867;
cipher_text[44] = `CIPHERTEXT_WIDTH'd15395717;
cipher_text[45] = `CIPHERTEXT_WIDTH'd10197904;
cipher_text[46] = `CIPHERTEXT_WIDTH'd14775933;
cipher_text[47] = `CIPHERTEXT_WIDTH'd2459182;
cipher_text[48] = `CIPHERTEXT_WIDTH'd2371464;
cipher_text[49] = `CIPHERTEXT_WIDTH'd360901;
cipher_text[50] = `CIPHERTEXT_WIDTH'd5790156;
cipher_text[51] = `CIPHERTEXT_WIDTH'd15659920;
cipher_text[52] = `CIPHERTEXT_WIDTH'd1390354;
cipher_text[53] = `CIPHERTEXT_WIDTH'd5987255;
cipher_text[54] = `CIPHERTEXT_WIDTH'd3829651;
cipher_text[55] = `CIPHERTEXT_WIDTH'd14490834;
cipher_text[56] = `CIPHERTEXT_WIDTH'd8144183;
cipher_text[57] = `CIPHERTEXT_WIDTH'd6250281;
cipher_text[58] = `CIPHERTEXT_WIDTH'd12816188;
cipher_text[59] = `CIPHERTEXT_WIDTH'd8254660;
cipher_text[60] = `CIPHERTEXT_WIDTH'd16252741;
cipher_text[61] = `CIPHERTEXT_WIDTH'd1271337;
cipher_text[62] = `CIPHERTEXT_WIDTH'd5970351;
cipher_text[63] = `CIPHERTEXT_WIDTH'd2548638;
cipher_text[64] = `CIPHERTEXT_WIDTH'd3391051;
cipher_text[65] = `CIPHERTEXT_WIDTH'd1541582;
cipher_text[66] = `CIPHERTEXT_WIDTH'd11967716;
cipher_text[67] = `CIPHERTEXT_WIDTH'd7954996;
cipher_text[68] = `CIPHERTEXT_WIDTH'd1787684;
cipher_text[69] = `CIPHERTEXT_WIDTH'd14067825;
cipher_text[70] = `CIPHERTEXT_WIDTH'd13278168;
cipher_text[71] = `CIPHERTEXT_WIDTH'd10878571;
cipher_text[72] = `CIPHERTEXT_WIDTH'd12043529;
cipher_text[73] = `CIPHERTEXT_WIDTH'd4933725;
cipher_text[74] = `CIPHERTEXT_WIDTH'd3102663;
cipher_text[75] = `CIPHERTEXT_WIDTH'd6666532;
cipher_text[76] = `CIPHERTEXT_WIDTH'd636683;
cipher_text[77] = `CIPHERTEXT_WIDTH'd2757868;
cipher_text[78] = `CIPHERTEXT_WIDTH'd1546180;
cipher_text[79] = `CIPHERTEXT_WIDTH'd12727579;
cipher_text[80] = `CIPHERTEXT_WIDTH'd3202912;
cipher_text[81] = `CIPHERTEXT_WIDTH'd12275544;
cipher_text[82] = `CIPHERTEXT_WIDTH'd1545388;
cipher_text[83] = `CIPHERTEXT_WIDTH'd8911806;
cipher_text[84] = `CIPHERTEXT_WIDTH'd4553534;
cipher_text[85] = `CIPHERTEXT_WIDTH'd12233508;
cipher_text[86] = `CIPHERTEXT_WIDTH'd14142931;
cipher_text[87] = `CIPHERTEXT_WIDTH'd16099527;
cipher_text[88] = `CIPHERTEXT_WIDTH'd8158973;
cipher_text[89] = `CIPHERTEXT_WIDTH'd14441151;
cipher_text[90] = `CIPHERTEXT_WIDTH'd7871513;
cipher_text[91] = `CIPHERTEXT_WIDTH'd15973872;
cipher_text[92] = `CIPHERTEXT_WIDTH'd10711522;
cipher_text[93] = `CIPHERTEXT_WIDTH'd2308491;
cipher_text[94] = `CIPHERTEXT_WIDTH'd2621706;
cipher_text[95] = `CIPHERTEXT_WIDTH'd6900965;
cipher_text[96] = `CIPHERTEXT_WIDTH'd6550437;
cipher_text[97] = `CIPHERTEXT_WIDTH'd15675495;
cipher_text[98] = `CIPHERTEXT_WIDTH'd12525757;
cipher_text[99] = `CIPHERTEXT_WIDTH'd16318036;
cipher_text[100] = `CIPHERTEXT_WIDTH'd11679560;
cipher_text[101] = `CIPHERTEXT_WIDTH'd4387625;
cipher_text[102] = `CIPHERTEXT_WIDTH'd12486051;
cipher_text[103] = `CIPHERTEXT_WIDTH'd12279568;
cipher_text[104] = `CIPHERTEXT_WIDTH'd8728776;
cipher_text[105] = `CIPHERTEXT_WIDTH'd10470959;
cipher_text[106] = `CIPHERTEXT_WIDTH'd8314586;
cipher_text[107] = `CIPHERTEXT_WIDTH'd1178083;
cipher_text[108] = `CIPHERTEXT_WIDTH'd13262923;
cipher_text[109] = `CIPHERTEXT_WIDTH'd1371527;
cipher_text[110] = `CIPHERTEXT_WIDTH'd256272;
cipher_text[111] = `CIPHERTEXT_WIDTH'd9979270;
cipher_text[112] = `CIPHERTEXT_WIDTH'd8127788;
cipher_text[113] = `CIPHERTEXT_WIDTH'd16290937;
cipher_text[114] = `CIPHERTEXT_WIDTH'd2860952;
cipher_text[115] = `CIPHERTEXT_WIDTH'd9197485;
cipher_text[116] = `CIPHERTEXT_WIDTH'd5836319;
cipher_text[117] = `CIPHERTEXT_WIDTH'd10917562;
cipher_text[118] = `CIPHERTEXT_WIDTH'd13337437;
cipher_text[119] = `CIPHERTEXT_WIDTH'd12374985;
cipher_text[120] = `CIPHERTEXT_WIDTH'd5530198;
cipher_text[121] = `CIPHERTEXT_WIDTH'd11293171;
cipher_text[122] = `CIPHERTEXT_WIDTH'd5373522;
cipher_text[123] = `CIPHERTEXT_WIDTH'd8388725;
cipher_text[124] = `CIPHERTEXT_WIDTH'd16485520;
cipher_text[125] = `CIPHERTEXT_WIDTH'd2677350;
cipher_text[126] = `CIPHERTEXT_WIDTH'd11730863;
cipher_text[127] = `CIPHERTEXT_WIDTH'd10163811;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 13;
cipher_text[0] = `CIPHERTEXT_WIDTH'd13244420;
cipher_text[1] = `CIPHERTEXT_WIDTH'd5897693;
cipher_text[2] = `CIPHERTEXT_WIDTH'd16492020;
cipher_text[3] = `CIPHERTEXT_WIDTH'd8522059;
cipher_text[4] = `CIPHERTEXT_WIDTH'd8132063;
cipher_text[5] = `CIPHERTEXT_WIDTH'd8316364;
cipher_text[6] = `CIPHERTEXT_WIDTH'd10418199;
cipher_text[7] = `CIPHERTEXT_WIDTH'd6071182;
cipher_text[8] = `CIPHERTEXT_WIDTH'd5934812;
cipher_text[9] = `CIPHERTEXT_WIDTH'd10423974;
cipher_text[10] = `CIPHERTEXT_WIDTH'd8059533;
cipher_text[11] = `CIPHERTEXT_WIDTH'd15866095;
cipher_text[12] = `CIPHERTEXT_WIDTH'd5505912;
cipher_text[13] = `CIPHERTEXT_WIDTH'd12534597;
cipher_text[14] = `CIPHERTEXT_WIDTH'd16267315;
cipher_text[15] = `CIPHERTEXT_WIDTH'd2551926;
cipher_text[16] = `CIPHERTEXT_WIDTH'd10971174;
cipher_text[17] = `CIPHERTEXT_WIDTH'd15533363;
cipher_text[18] = `CIPHERTEXT_WIDTH'd6567060;
cipher_text[19] = `CIPHERTEXT_WIDTH'd14339001;
cipher_text[20] = `CIPHERTEXT_WIDTH'd14254862;
cipher_text[21] = `CIPHERTEXT_WIDTH'd9210297;
cipher_text[22] = `CIPHERTEXT_WIDTH'd13903516;
cipher_text[23] = `CIPHERTEXT_WIDTH'd6384514;
cipher_text[24] = `CIPHERTEXT_WIDTH'd16012539;
cipher_text[25] = `CIPHERTEXT_WIDTH'd9590018;
cipher_text[26] = `CIPHERTEXT_WIDTH'd9436168;
cipher_text[27] = `CIPHERTEXT_WIDTH'd12561402;
cipher_text[28] = `CIPHERTEXT_WIDTH'd16107039;
cipher_text[29] = `CIPHERTEXT_WIDTH'd9210802;
cipher_text[30] = `CIPHERTEXT_WIDTH'd8866860;
cipher_text[31] = `CIPHERTEXT_WIDTH'd15752838;
cipher_text[32] = `CIPHERTEXT_WIDTH'd8113233;
cipher_text[33] = `CIPHERTEXT_WIDTH'd5574666;
cipher_text[34] = `CIPHERTEXT_WIDTH'd13053604;
cipher_text[35] = `CIPHERTEXT_WIDTH'd2374094;
cipher_text[36] = `CIPHERTEXT_WIDTH'd10049527;
cipher_text[37] = `CIPHERTEXT_WIDTH'd2539974;
cipher_text[38] = `CIPHERTEXT_WIDTH'd10531372;
cipher_text[39] = `CIPHERTEXT_WIDTH'd2975473;
cipher_text[40] = `CIPHERTEXT_WIDTH'd14128809;
cipher_text[41] = `CIPHERTEXT_WIDTH'd10651179;
cipher_text[42] = `CIPHERTEXT_WIDTH'd10422345;
cipher_text[43] = `CIPHERTEXT_WIDTH'd8869085;
cipher_text[44] = `CIPHERTEXT_WIDTH'd15751560;
cipher_text[45] = `CIPHERTEXT_WIDTH'd3496490;
cipher_text[46] = `CIPHERTEXT_WIDTH'd541787;
cipher_text[47] = `CIPHERTEXT_WIDTH'd766875;
cipher_text[48] = `CIPHERTEXT_WIDTH'd13399225;
cipher_text[49] = `CIPHERTEXT_WIDTH'd10832082;
cipher_text[50] = `CIPHERTEXT_WIDTH'd6048676;
cipher_text[51] = `CIPHERTEXT_WIDTH'd5612380;
cipher_text[52] = `CIPHERTEXT_WIDTH'd5340631;
cipher_text[53] = `CIPHERTEXT_WIDTH'd15501823;
cipher_text[54] = `CIPHERTEXT_WIDTH'd12386133;
cipher_text[55] = `CIPHERTEXT_WIDTH'd4892829;
cipher_text[56] = `CIPHERTEXT_WIDTH'd1717564;
cipher_text[57] = `CIPHERTEXT_WIDTH'd1018173;
cipher_text[58] = `CIPHERTEXT_WIDTH'd8698730;
cipher_text[59] = `CIPHERTEXT_WIDTH'd16231162;
cipher_text[60] = `CIPHERTEXT_WIDTH'd12975641;
cipher_text[61] = `CIPHERTEXT_WIDTH'd16108728;
cipher_text[62] = `CIPHERTEXT_WIDTH'd14690464;
cipher_text[63] = `CIPHERTEXT_WIDTH'd15673831;
cipher_text[64] = `CIPHERTEXT_WIDTH'd10551308;
cipher_text[65] = `CIPHERTEXT_WIDTH'd6898904;
cipher_text[66] = `CIPHERTEXT_WIDTH'd1699139;
cipher_text[67] = `CIPHERTEXT_WIDTH'd12554371;
cipher_text[68] = `CIPHERTEXT_WIDTH'd5308666;
cipher_text[69] = `CIPHERTEXT_WIDTH'd8095091;
cipher_text[70] = `CIPHERTEXT_WIDTH'd1991091;
cipher_text[71] = `CIPHERTEXT_WIDTH'd6721744;
cipher_text[72] = `CIPHERTEXT_WIDTH'd10981716;
cipher_text[73] = `CIPHERTEXT_WIDTH'd15807917;
cipher_text[74] = `CIPHERTEXT_WIDTH'd5143300;
cipher_text[75] = `CIPHERTEXT_WIDTH'd1281340;
cipher_text[76] = `CIPHERTEXT_WIDTH'd4467206;
cipher_text[77] = `CIPHERTEXT_WIDTH'd1767427;
cipher_text[78] = `CIPHERTEXT_WIDTH'd9018811;
cipher_text[79] = `CIPHERTEXT_WIDTH'd2966678;
cipher_text[80] = `CIPHERTEXT_WIDTH'd16697240;
cipher_text[81] = `CIPHERTEXT_WIDTH'd10779366;
cipher_text[82] = `CIPHERTEXT_WIDTH'd12620357;
cipher_text[83] = `CIPHERTEXT_WIDTH'd1897807;
cipher_text[84] = `CIPHERTEXT_WIDTH'd11648534;
cipher_text[85] = `CIPHERTEXT_WIDTH'd4776603;
cipher_text[86] = `CIPHERTEXT_WIDTH'd14303510;
cipher_text[87] = `CIPHERTEXT_WIDTH'd16069899;
cipher_text[88] = `CIPHERTEXT_WIDTH'd4413167;
cipher_text[89] = `CIPHERTEXT_WIDTH'd6683364;
cipher_text[90] = `CIPHERTEXT_WIDTH'd15397816;
cipher_text[91] = `CIPHERTEXT_WIDTH'd3309833;
cipher_text[92] = `CIPHERTEXT_WIDTH'd5856834;
cipher_text[93] = `CIPHERTEXT_WIDTH'd11967605;
cipher_text[94] = `CIPHERTEXT_WIDTH'd6441444;
cipher_text[95] = `CIPHERTEXT_WIDTH'd15541036;
cipher_text[96] = `CIPHERTEXT_WIDTH'd4010395;
cipher_text[97] = `CIPHERTEXT_WIDTH'd12074559;
cipher_text[98] = `CIPHERTEXT_WIDTH'd5173018;
cipher_text[99] = `CIPHERTEXT_WIDTH'd3546559;
cipher_text[100] = `CIPHERTEXT_WIDTH'd1925250;
cipher_text[101] = `CIPHERTEXT_WIDTH'd15196890;
cipher_text[102] = `CIPHERTEXT_WIDTH'd1338840;
cipher_text[103] = `CIPHERTEXT_WIDTH'd5659063;
cipher_text[104] = `CIPHERTEXT_WIDTH'd12707098;
cipher_text[105] = `CIPHERTEXT_WIDTH'd3538555;
cipher_text[106] = `CIPHERTEXT_WIDTH'd1407436;
cipher_text[107] = `CIPHERTEXT_WIDTH'd4966515;
cipher_text[108] = `CIPHERTEXT_WIDTH'd13415997;
cipher_text[109] = `CIPHERTEXT_WIDTH'd163526;
cipher_text[110] = `CIPHERTEXT_WIDTH'd9311802;
cipher_text[111] = `CIPHERTEXT_WIDTH'd10442008;
cipher_text[112] = `CIPHERTEXT_WIDTH'd12004606;
cipher_text[113] = `CIPHERTEXT_WIDTH'd12509496;
cipher_text[114] = `CIPHERTEXT_WIDTH'd13013654;
cipher_text[115] = `CIPHERTEXT_WIDTH'd9359322;
cipher_text[116] = `CIPHERTEXT_WIDTH'd8409786;
cipher_text[117] = `CIPHERTEXT_WIDTH'd1986218;
cipher_text[118] = `CIPHERTEXT_WIDTH'd9077559;
cipher_text[119] = `CIPHERTEXT_WIDTH'd10944071;
cipher_text[120] = `CIPHERTEXT_WIDTH'd5948802;
cipher_text[121] = `CIPHERTEXT_WIDTH'd522963;
cipher_text[122] = `CIPHERTEXT_WIDTH'd8858265;
cipher_text[123] = `CIPHERTEXT_WIDTH'd4206188;
cipher_text[124] = `CIPHERTEXT_WIDTH'd9018963;
cipher_text[125] = `CIPHERTEXT_WIDTH'd11154892;
cipher_text[126] = `CIPHERTEXT_WIDTH'd2821252;
cipher_text[127] = `CIPHERTEXT_WIDTH'd13501864;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 14;
cipher_text[0] = `CIPHERTEXT_WIDTH'd13333932;
cipher_text[1] = `CIPHERTEXT_WIDTH'd3561209;
cipher_text[2] = `CIPHERTEXT_WIDTH'd9815128;
cipher_text[3] = `CIPHERTEXT_WIDTH'd16723164;
cipher_text[4] = `CIPHERTEXT_WIDTH'd12260520;
cipher_text[5] = `CIPHERTEXT_WIDTH'd8838427;
cipher_text[6] = `CIPHERTEXT_WIDTH'd8360253;
cipher_text[7] = `CIPHERTEXT_WIDTH'd3761243;
cipher_text[8] = `CIPHERTEXT_WIDTH'd3926445;
cipher_text[9] = `CIPHERTEXT_WIDTH'd7628192;
cipher_text[10] = `CIPHERTEXT_WIDTH'd15632690;
cipher_text[11] = `CIPHERTEXT_WIDTH'd3701110;
cipher_text[12] = `CIPHERTEXT_WIDTH'd16475220;
cipher_text[13] = `CIPHERTEXT_WIDTH'd2941959;
cipher_text[14] = `CIPHERTEXT_WIDTH'd12548415;
cipher_text[15] = `CIPHERTEXT_WIDTH'd10926701;
cipher_text[16] = `CIPHERTEXT_WIDTH'd11667399;
cipher_text[17] = `CIPHERTEXT_WIDTH'd4728183;
cipher_text[18] = `CIPHERTEXT_WIDTH'd979834;
cipher_text[19] = `CIPHERTEXT_WIDTH'd15779752;
cipher_text[20] = `CIPHERTEXT_WIDTH'd3302487;
cipher_text[21] = `CIPHERTEXT_WIDTH'd3329223;
cipher_text[22] = `CIPHERTEXT_WIDTH'd932296;
cipher_text[23] = `CIPHERTEXT_WIDTH'd9380692;
cipher_text[24] = `CIPHERTEXT_WIDTH'd16036709;
cipher_text[25] = `CIPHERTEXT_WIDTH'd524053;
cipher_text[26] = `CIPHERTEXT_WIDTH'd479568;
cipher_text[27] = `CIPHERTEXT_WIDTH'd865212;
cipher_text[28] = `CIPHERTEXT_WIDTH'd16064068;
cipher_text[29] = `CIPHERTEXT_WIDTH'd16579537;
cipher_text[30] = `CIPHERTEXT_WIDTH'd2069921;
cipher_text[31] = `CIPHERTEXT_WIDTH'd11404155;
cipher_text[32] = `CIPHERTEXT_WIDTH'd9350535;
cipher_text[33] = `CIPHERTEXT_WIDTH'd15982788;
cipher_text[34] = `CIPHERTEXT_WIDTH'd3553954;
cipher_text[35] = `CIPHERTEXT_WIDTH'd9832247;
cipher_text[36] = `CIPHERTEXT_WIDTH'd11537850;
cipher_text[37] = `CIPHERTEXT_WIDTH'd172309;
cipher_text[38] = `CIPHERTEXT_WIDTH'd9193361;
cipher_text[39] = `CIPHERTEXT_WIDTH'd5437993;
cipher_text[40] = `CIPHERTEXT_WIDTH'd15405977;
cipher_text[41] = `CIPHERTEXT_WIDTH'd667621;
cipher_text[42] = `CIPHERTEXT_WIDTH'd6313142;
cipher_text[43] = `CIPHERTEXT_WIDTH'd12640240;
cipher_text[44] = `CIPHERTEXT_WIDTH'd11544757;
cipher_text[45] = `CIPHERTEXT_WIDTH'd10876118;
cipher_text[46] = `CIPHERTEXT_WIDTH'd3083992;
cipher_text[47] = `CIPHERTEXT_WIDTH'd8827993;
cipher_text[48] = `CIPHERTEXT_WIDTH'd5922290;
cipher_text[49] = `CIPHERTEXT_WIDTH'd7316996;
cipher_text[50] = `CIPHERTEXT_WIDTH'd16303837;
cipher_text[51] = `CIPHERTEXT_WIDTH'd10696090;
cipher_text[52] = `CIPHERTEXT_WIDTH'd11854199;
cipher_text[53] = `CIPHERTEXT_WIDTH'd8264035;
cipher_text[54] = `CIPHERTEXT_WIDTH'd16438638;
cipher_text[55] = `CIPHERTEXT_WIDTH'd11711901;
cipher_text[56] = `CIPHERTEXT_WIDTH'd2700982;
cipher_text[57] = `CIPHERTEXT_WIDTH'd9431876;
cipher_text[58] = `CIPHERTEXT_WIDTH'd5447689;
cipher_text[59] = `CIPHERTEXT_WIDTH'd15060865;
cipher_text[60] = `CIPHERTEXT_WIDTH'd1628742;
cipher_text[61] = `CIPHERTEXT_WIDTH'd359747;
cipher_text[62] = `CIPHERTEXT_WIDTH'd1990750;
cipher_text[63] = `CIPHERTEXT_WIDTH'd4912554;
cipher_text[64] = `CIPHERTEXT_WIDTH'd9250331;
cipher_text[65] = `CIPHERTEXT_WIDTH'd6291799;
cipher_text[66] = `CIPHERTEXT_WIDTH'd12485356;
cipher_text[67] = `CIPHERTEXT_WIDTH'd2158601;
cipher_text[68] = `CIPHERTEXT_WIDTH'd14565330;
cipher_text[69] = `CIPHERTEXT_WIDTH'd11067280;
cipher_text[70] = `CIPHERTEXT_WIDTH'd9183684;
cipher_text[71] = `CIPHERTEXT_WIDTH'd12742167;
cipher_text[72] = `CIPHERTEXT_WIDTH'd13021414;
cipher_text[73] = `CIPHERTEXT_WIDTH'd12520505;
cipher_text[74] = `CIPHERTEXT_WIDTH'd5405600;
cipher_text[75] = `CIPHERTEXT_WIDTH'd11032022;
cipher_text[76] = `CIPHERTEXT_WIDTH'd8600157;
cipher_text[77] = `CIPHERTEXT_WIDTH'd8549406;
cipher_text[78] = `CIPHERTEXT_WIDTH'd7892988;
cipher_text[79] = `CIPHERTEXT_WIDTH'd10060267;
cipher_text[80] = `CIPHERTEXT_WIDTH'd10559828;
cipher_text[81] = `CIPHERTEXT_WIDTH'd12760178;
cipher_text[82] = `CIPHERTEXT_WIDTH'd4361031;
cipher_text[83] = `CIPHERTEXT_WIDTH'd663213;
cipher_text[84] = `CIPHERTEXT_WIDTH'd2256099;
cipher_text[85] = `CIPHERTEXT_WIDTH'd13568419;
cipher_text[86] = `CIPHERTEXT_WIDTH'd12092063;
cipher_text[87] = `CIPHERTEXT_WIDTH'd5156938;
cipher_text[88] = `CIPHERTEXT_WIDTH'd11863428;
cipher_text[89] = `CIPHERTEXT_WIDTH'd10746454;
cipher_text[90] = `CIPHERTEXT_WIDTH'd14086651;
cipher_text[91] = `CIPHERTEXT_WIDTH'd603196;
cipher_text[92] = `CIPHERTEXT_WIDTH'd12226025;
cipher_text[93] = `CIPHERTEXT_WIDTH'd3672981;
cipher_text[94] = `CIPHERTEXT_WIDTH'd500298;
cipher_text[95] = `CIPHERTEXT_WIDTH'd14896271;
cipher_text[96] = `CIPHERTEXT_WIDTH'd10287639;
cipher_text[97] = `CIPHERTEXT_WIDTH'd9498689;
cipher_text[98] = `CIPHERTEXT_WIDTH'd10285130;
cipher_text[99] = `CIPHERTEXT_WIDTH'd10047584;
cipher_text[100] = `CIPHERTEXT_WIDTH'd2360662;
cipher_text[101] = `CIPHERTEXT_WIDTH'd3847761;
cipher_text[102] = `CIPHERTEXT_WIDTH'd6254178;
cipher_text[103] = `CIPHERTEXT_WIDTH'd6526237;
cipher_text[104] = `CIPHERTEXT_WIDTH'd15174046;
cipher_text[105] = `CIPHERTEXT_WIDTH'd172857;
cipher_text[106] = `CIPHERTEXT_WIDTH'd811432;
cipher_text[107] = `CIPHERTEXT_WIDTH'd15013268;
cipher_text[108] = `CIPHERTEXT_WIDTH'd4437292;
cipher_text[109] = `CIPHERTEXT_WIDTH'd11290858;
cipher_text[110] = `CIPHERTEXT_WIDTH'd12076353;
cipher_text[111] = `CIPHERTEXT_WIDTH'd4328605;
cipher_text[112] = `CIPHERTEXT_WIDTH'd8871740;
cipher_text[113] = `CIPHERTEXT_WIDTH'd8793875;
cipher_text[114] = `CIPHERTEXT_WIDTH'd1607326;
cipher_text[115] = `CIPHERTEXT_WIDTH'd6049940;
cipher_text[116] = `CIPHERTEXT_WIDTH'd1037564;
cipher_text[117] = `CIPHERTEXT_WIDTH'd12109220;
cipher_text[118] = `CIPHERTEXT_WIDTH'd12853112;
cipher_text[119] = `CIPHERTEXT_WIDTH'd4433207;
cipher_text[120] = `CIPHERTEXT_WIDTH'd4031904;
cipher_text[121] = `CIPHERTEXT_WIDTH'd2929654;
cipher_text[122] = `CIPHERTEXT_WIDTH'd11274638;
cipher_text[123] = `CIPHERTEXT_WIDTH'd1850033;
cipher_text[124] = `CIPHERTEXT_WIDTH'd5009755;
cipher_text[125] = `CIPHERTEXT_WIDTH'd14453475;
cipher_text[126] = `CIPHERTEXT_WIDTH'd8187752;
cipher_text[127] = `CIPHERTEXT_WIDTH'd11628871;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 15;
cipher_text[0] = `CIPHERTEXT_WIDTH'd13760424;
cipher_text[1] = `CIPHERTEXT_WIDTH'd3652529;
cipher_text[2] = `CIPHERTEXT_WIDTH'd11397337;
cipher_text[3] = `CIPHERTEXT_WIDTH'd4312539;
cipher_text[4] = `CIPHERTEXT_WIDTH'd7854533;
cipher_text[5] = `CIPHERTEXT_WIDTH'd14482580;
cipher_text[6] = `CIPHERTEXT_WIDTH'd3362018;
cipher_text[7] = `CIPHERTEXT_WIDTH'd11924900;
cipher_text[8] = `CIPHERTEXT_WIDTH'd10707003;
cipher_text[9] = `CIPHERTEXT_WIDTH'd6633090;
cipher_text[10] = `CIPHERTEXT_WIDTH'd10005338;
cipher_text[11] = `CIPHERTEXT_WIDTH'd16157048;
cipher_text[12] = `CIPHERTEXT_WIDTH'd15428834;
cipher_text[13] = `CIPHERTEXT_WIDTH'd1873170;
cipher_text[14] = `CIPHERTEXT_WIDTH'd2298612;
cipher_text[15] = `CIPHERTEXT_WIDTH'd10964987;
cipher_text[16] = `CIPHERTEXT_WIDTH'd6972126;
cipher_text[17] = `CIPHERTEXT_WIDTH'd15806658;
cipher_text[18] = `CIPHERTEXT_WIDTH'd1554768;
cipher_text[19] = `CIPHERTEXT_WIDTH'd12350235;
cipher_text[20] = `CIPHERTEXT_WIDTH'd11717735;
cipher_text[21] = `CIPHERTEXT_WIDTH'd11095799;
cipher_text[22] = `CIPHERTEXT_WIDTH'd10520105;
cipher_text[23] = `CIPHERTEXT_WIDTH'd1742616;
cipher_text[24] = `CIPHERTEXT_WIDTH'd4011777;
cipher_text[25] = `CIPHERTEXT_WIDTH'd6659329;
cipher_text[26] = `CIPHERTEXT_WIDTH'd3554121;
cipher_text[27] = `CIPHERTEXT_WIDTH'd13415450;
cipher_text[28] = `CIPHERTEXT_WIDTH'd13449574;
cipher_text[29] = `CIPHERTEXT_WIDTH'd8705387;
cipher_text[30] = `CIPHERTEXT_WIDTH'd2931628;
cipher_text[31] = `CIPHERTEXT_WIDTH'd16507740;
cipher_text[32] = `CIPHERTEXT_WIDTH'd3624489;
cipher_text[33] = `CIPHERTEXT_WIDTH'd9183466;
cipher_text[34] = `CIPHERTEXT_WIDTH'd1234611;
cipher_text[35] = `CIPHERTEXT_WIDTH'd11769229;
cipher_text[36] = `CIPHERTEXT_WIDTH'd4024795;
cipher_text[37] = `CIPHERTEXT_WIDTH'd1831326;
cipher_text[38] = `CIPHERTEXT_WIDTH'd8603570;
cipher_text[39] = `CIPHERTEXT_WIDTH'd15465455;
cipher_text[40] = `CIPHERTEXT_WIDTH'd6293491;
cipher_text[41] = `CIPHERTEXT_WIDTH'd12490875;
cipher_text[42] = `CIPHERTEXT_WIDTH'd4064878;
cipher_text[43] = `CIPHERTEXT_WIDTH'd13966083;
cipher_text[44] = `CIPHERTEXT_WIDTH'd8651697;
cipher_text[45] = `CIPHERTEXT_WIDTH'd12644514;
cipher_text[46] = `CIPHERTEXT_WIDTH'd6877851;
cipher_text[47] = `CIPHERTEXT_WIDTH'd15430312;
cipher_text[48] = `CIPHERTEXT_WIDTH'd4223188;
cipher_text[49] = `CIPHERTEXT_WIDTH'd10277907;
cipher_text[50] = `CIPHERTEXT_WIDTH'd7088544;
cipher_text[51] = `CIPHERTEXT_WIDTH'd1301325;
cipher_text[52] = `CIPHERTEXT_WIDTH'd8644678;
cipher_text[53] = `CIPHERTEXT_WIDTH'd3306822;
cipher_text[54] = `CIPHERTEXT_WIDTH'd13915169;
cipher_text[55] = `CIPHERTEXT_WIDTH'd10394055;
cipher_text[56] = `CIPHERTEXT_WIDTH'd5726392;
cipher_text[57] = `CIPHERTEXT_WIDTH'd9327658;
cipher_text[58] = `CIPHERTEXT_WIDTH'd1976176;
cipher_text[59] = `CIPHERTEXT_WIDTH'd11779338;
cipher_text[60] = `CIPHERTEXT_WIDTH'd8062260;
cipher_text[61] = `CIPHERTEXT_WIDTH'd7592747;
cipher_text[62] = `CIPHERTEXT_WIDTH'd2528022;
cipher_text[63] = `CIPHERTEXT_WIDTH'd11987315;
cipher_text[64] = `CIPHERTEXT_WIDTH'd11372766;
cipher_text[65] = `CIPHERTEXT_WIDTH'd2269993;
cipher_text[66] = `CIPHERTEXT_WIDTH'd2403880;
cipher_text[67] = `CIPHERTEXT_WIDTH'd8628507;
cipher_text[68] = `CIPHERTEXT_WIDTH'd937435;
cipher_text[69] = `CIPHERTEXT_WIDTH'd7546707;
cipher_text[70] = `CIPHERTEXT_WIDTH'd4091632;
cipher_text[71] = `CIPHERTEXT_WIDTH'd14377045;
cipher_text[72] = `CIPHERTEXT_WIDTH'd15873276;
cipher_text[73] = `CIPHERTEXT_WIDTH'd16741909;
cipher_text[74] = `CIPHERTEXT_WIDTH'd12979120;
cipher_text[75] = `CIPHERTEXT_WIDTH'd14639373;
cipher_text[76] = `CIPHERTEXT_WIDTH'd11714427;
cipher_text[77] = `CIPHERTEXT_WIDTH'd499729;
cipher_text[78] = `CIPHERTEXT_WIDTH'd13118655;
cipher_text[79] = `CIPHERTEXT_WIDTH'd13004196;
cipher_text[80] = `CIPHERTEXT_WIDTH'd1460705;
cipher_text[81] = `CIPHERTEXT_WIDTH'd8773160;
cipher_text[82] = `CIPHERTEXT_WIDTH'd4218401;
cipher_text[83] = `CIPHERTEXT_WIDTH'd12273687;
cipher_text[84] = `CIPHERTEXT_WIDTH'd4907382;
cipher_text[85] = `CIPHERTEXT_WIDTH'd13918458;
cipher_text[86] = `CIPHERTEXT_WIDTH'd6143997;
cipher_text[87] = `CIPHERTEXT_WIDTH'd1105845;
cipher_text[88] = `CIPHERTEXT_WIDTH'd14433792;
cipher_text[89] = `CIPHERTEXT_WIDTH'd12110871;
cipher_text[90] = `CIPHERTEXT_WIDTH'd12661029;
cipher_text[91] = `CIPHERTEXT_WIDTH'd944526;
cipher_text[92] = `CIPHERTEXT_WIDTH'd15714618;
cipher_text[93] = `CIPHERTEXT_WIDTH'd1119634;
cipher_text[94] = `CIPHERTEXT_WIDTH'd12312029;
cipher_text[95] = `CIPHERTEXT_WIDTH'd7145775;
cipher_text[96] = `CIPHERTEXT_WIDTH'd8762677;
cipher_text[97] = `CIPHERTEXT_WIDTH'd3670651;
cipher_text[98] = `CIPHERTEXT_WIDTH'd5546990;
cipher_text[99] = `CIPHERTEXT_WIDTH'd5687028;
cipher_text[100] = `CIPHERTEXT_WIDTH'd10286269;
cipher_text[101] = `CIPHERTEXT_WIDTH'd13402767;
cipher_text[102] = `CIPHERTEXT_WIDTH'd12309327;
cipher_text[103] = `CIPHERTEXT_WIDTH'd15783656;
cipher_text[104] = `CIPHERTEXT_WIDTH'd14950504;
cipher_text[105] = `CIPHERTEXT_WIDTH'd7368132;
cipher_text[106] = `CIPHERTEXT_WIDTH'd1009364;
cipher_text[107] = `CIPHERTEXT_WIDTH'd107703;
cipher_text[108] = `CIPHERTEXT_WIDTH'd5809136;
cipher_text[109] = `CIPHERTEXT_WIDTH'd4447916;
cipher_text[110] = `CIPHERTEXT_WIDTH'd2689628;
cipher_text[111] = `CIPHERTEXT_WIDTH'd8600127;
cipher_text[112] = `CIPHERTEXT_WIDTH'd14315653;
cipher_text[113] = `CIPHERTEXT_WIDTH'd7311702;
cipher_text[114] = `CIPHERTEXT_WIDTH'd3480457;
cipher_text[115] = `CIPHERTEXT_WIDTH'd12194572;
cipher_text[116] = `CIPHERTEXT_WIDTH'd668606;
cipher_text[117] = `CIPHERTEXT_WIDTH'd9402177;
cipher_text[118] = `CIPHERTEXT_WIDTH'd6553222;
cipher_text[119] = `CIPHERTEXT_WIDTH'd15076566;
cipher_text[120] = `CIPHERTEXT_WIDTH'd16260108;
cipher_text[121] = `CIPHERTEXT_WIDTH'd8722197;
cipher_text[122] = `CIPHERTEXT_WIDTH'd15918756;
cipher_text[123] = `CIPHERTEXT_WIDTH'd2015238;
cipher_text[124] = `CIPHERTEXT_WIDTH'd3932385;
cipher_text[125] = `CIPHERTEXT_WIDTH'd8649791;
cipher_text[126] = `CIPHERTEXT_WIDTH'd2899755;
cipher_text[127] = `CIPHERTEXT_WIDTH'd11168250;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 16;
cipher_text[0] = `CIPHERTEXT_WIDTH'd9857588;
cipher_text[1] = `CIPHERTEXT_WIDTH'd6350545;
cipher_text[2] = `CIPHERTEXT_WIDTH'd10618476;
cipher_text[3] = `CIPHERTEXT_WIDTH'd13591628;
cipher_text[4] = `CIPHERTEXT_WIDTH'd6971727;
cipher_text[5] = `CIPHERTEXT_WIDTH'd7575062;
cipher_text[6] = `CIPHERTEXT_WIDTH'd278348;
cipher_text[7] = `CIPHERTEXT_WIDTH'd7824360;
cipher_text[8] = `CIPHERTEXT_WIDTH'd16045864;
cipher_text[9] = `CIPHERTEXT_WIDTH'd5713501;
cipher_text[10] = `CIPHERTEXT_WIDTH'd14948352;
cipher_text[11] = `CIPHERTEXT_WIDTH'd6687868;
cipher_text[12] = `CIPHERTEXT_WIDTH'd4427804;
cipher_text[13] = `CIPHERTEXT_WIDTH'd14521620;
cipher_text[14] = `CIPHERTEXT_WIDTH'd10320683;
cipher_text[15] = `CIPHERTEXT_WIDTH'd16344698;
cipher_text[16] = `CIPHERTEXT_WIDTH'd3250311;
cipher_text[17] = `CIPHERTEXT_WIDTH'd5098399;
cipher_text[18] = `CIPHERTEXT_WIDTH'd5743322;
cipher_text[19] = `CIPHERTEXT_WIDTH'd9560035;
cipher_text[20] = `CIPHERTEXT_WIDTH'd9160837;
cipher_text[21] = `CIPHERTEXT_WIDTH'd11237383;
cipher_text[22] = `CIPHERTEXT_WIDTH'd7138279;
cipher_text[23] = `CIPHERTEXT_WIDTH'd5900466;
cipher_text[24] = `CIPHERTEXT_WIDTH'd641511;
cipher_text[25] = `CIPHERTEXT_WIDTH'd11970323;
cipher_text[26] = `CIPHERTEXT_WIDTH'd4265245;
cipher_text[27] = `CIPHERTEXT_WIDTH'd344421;
cipher_text[28] = `CIPHERTEXT_WIDTH'd6971394;
cipher_text[29] = `CIPHERTEXT_WIDTH'd6718666;
cipher_text[30] = `CIPHERTEXT_WIDTH'd12774439;
cipher_text[31] = `CIPHERTEXT_WIDTH'd12384185;
cipher_text[32] = `CIPHERTEXT_WIDTH'd10750351;
cipher_text[33] = `CIPHERTEXT_WIDTH'd6873367;
cipher_text[34] = `CIPHERTEXT_WIDTH'd5655417;
cipher_text[35] = `CIPHERTEXT_WIDTH'd14649916;
cipher_text[36] = `CIPHERTEXT_WIDTH'd8992061;
cipher_text[37] = `CIPHERTEXT_WIDTH'd16776919;
cipher_text[38] = `CIPHERTEXT_WIDTH'd9257523;
cipher_text[39] = `CIPHERTEXT_WIDTH'd198258;
cipher_text[40] = `CIPHERTEXT_WIDTH'd15885180;
cipher_text[41] = `CIPHERTEXT_WIDTH'd1268894;
cipher_text[42] = `CIPHERTEXT_WIDTH'd13334349;
cipher_text[43] = `CIPHERTEXT_WIDTH'd6901526;
cipher_text[44] = `CIPHERTEXT_WIDTH'd12178119;
cipher_text[45] = `CIPHERTEXT_WIDTH'd16277625;
cipher_text[46] = `CIPHERTEXT_WIDTH'd1177351;
cipher_text[47] = `CIPHERTEXT_WIDTH'd9873112;
cipher_text[48] = `CIPHERTEXT_WIDTH'd11509362;
cipher_text[49] = `CIPHERTEXT_WIDTH'd9863615;
cipher_text[50] = `CIPHERTEXT_WIDTH'd4081154;
cipher_text[51] = `CIPHERTEXT_WIDTH'd5035920;
cipher_text[52] = `CIPHERTEXT_WIDTH'd2670314;
cipher_text[53] = `CIPHERTEXT_WIDTH'd15138151;
cipher_text[54] = `CIPHERTEXT_WIDTH'd14514878;
cipher_text[55] = `CIPHERTEXT_WIDTH'd11332944;
cipher_text[56] = `CIPHERTEXT_WIDTH'd9615804;
cipher_text[57] = `CIPHERTEXT_WIDTH'd7236723;
cipher_text[58] = `CIPHERTEXT_WIDTH'd2175319;
cipher_text[59] = `CIPHERTEXT_WIDTH'd2483800;
cipher_text[60] = `CIPHERTEXT_WIDTH'd8564470;
cipher_text[61] = `CIPHERTEXT_WIDTH'd14701988;
cipher_text[62] = `CIPHERTEXT_WIDTH'd9702170;
cipher_text[63] = `CIPHERTEXT_WIDTH'd4610254;
cipher_text[64] = `CIPHERTEXT_WIDTH'd13197243;
cipher_text[65] = `CIPHERTEXT_WIDTH'd4599597;
cipher_text[66] = `CIPHERTEXT_WIDTH'd6609452;
cipher_text[67] = `CIPHERTEXT_WIDTH'd1790469;
cipher_text[68] = `CIPHERTEXT_WIDTH'd8719607;
cipher_text[69] = `CIPHERTEXT_WIDTH'd13390555;
cipher_text[70] = `CIPHERTEXT_WIDTH'd16613906;
cipher_text[71] = `CIPHERTEXT_WIDTH'd3815275;
cipher_text[72] = `CIPHERTEXT_WIDTH'd491731;
cipher_text[73] = `CIPHERTEXT_WIDTH'd11305557;
cipher_text[74] = `CIPHERTEXT_WIDTH'd7754060;
cipher_text[75] = `CIPHERTEXT_WIDTH'd5446436;
cipher_text[76] = `CIPHERTEXT_WIDTH'd10002519;
cipher_text[77] = `CIPHERTEXT_WIDTH'd5337564;
cipher_text[78] = `CIPHERTEXT_WIDTH'd2492713;
cipher_text[79] = `CIPHERTEXT_WIDTH'd13016485;
cipher_text[80] = `CIPHERTEXT_WIDTH'd3849016;
cipher_text[81] = `CIPHERTEXT_WIDTH'd4579332;
cipher_text[82] = `CIPHERTEXT_WIDTH'd2351190;
cipher_text[83] = `CIPHERTEXT_WIDTH'd15703902;
cipher_text[84] = `CIPHERTEXT_WIDTH'd2284151;
cipher_text[85] = `CIPHERTEXT_WIDTH'd12906273;
cipher_text[86] = `CIPHERTEXT_WIDTH'd5541822;
cipher_text[87] = `CIPHERTEXT_WIDTH'd4951667;
cipher_text[88] = `CIPHERTEXT_WIDTH'd6482429;
cipher_text[89] = `CIPHERTEXT_WIDTH'd5948365;
cipher_text[90] = `CIPHERTEXT_WIDTH'd5022031;
cipher_text[91] = `CIPHERTEXT_WIDTH'd6971797;
cipher_text[92] = `CIPHERTEXT_WIDTH'd2666607;
cipher_text[93] = `CIPHERTEXT_WIDTH'd9399795;
cipher_text[94] = `CIPHERTEXT_WIDTH'd11620992;
cipher_text[95] = `CIPHERTEXT_WIDTH'd7117310;
cipher_text[96] = `CIPHERTEXT_WIDTH'd11158637;
cipher_text[97] = `CIPHERTEXT_WIDTH'd4168037;
cipher_text[98] = `CIPHERTEXT_WIDTH'd496166;
cipher_text[99] = `CIPHERTEXT_WIDTH'd14088291;
cipher_text[100] = `CIPHERTEXT_WIDTH'd212978;
cipher_text[101] = `CIPHERTEXT_WIDTH'd13669538;
cipher_text[102] = `CIPHERTEXT_WIDTH'd738637;
cipher_text[103] = `CIPHERTEXT_WIDTH'd10700943;
cipher_text[104] = `CIPHERTEXT_WIDTH'd10075324;
cipher_text[105] = `CIPHERTEXT_WIDTH'd2511928;
cipher_text[106] = `CIPHERTEXT_WIDTH'd3110540;
cipher_text[107] = `CIPHERTEXT_WIDTH'd12289163;
cipher_text[108] = `CIPHERTEXT_WIDTH'd11005253;
cipher_text[109] = `CIPHERTEXT_WIDTH'd11881674;
cipher_text[110] = `CIPHERTEXT_WIDTH'd10021396;
cipher_text[111] = `CIPHERTEXT_WIDTH'd10545689;
cipher_text[112] = `CIPHERTEXT_WIDTH'd8188136;
cipher_text[113] = `CIPHERTEXT_WIDTH'd7084847;
cipher_text[114] = `CIPHERTEXT_WIDTH'd6454674;
cipher_text[115] = `CIPHERTEXT_WIDTH'd11432879;
cipher_text[116] = `CIPHERTEXT_WIDTH'd7857433;
cipher_text[117] = `CIPHERTEXT_WIDTH'd694787;
cipher_text[118] = `CIPHERTEXT_WIDTH'd12897602;
cipher_text[119] = `CIPHERTEXT_WIDTH'd5510642;
cipher_text[120] = `CIPHERTEXT_WIDTH'd6245184;
cipher_text[121] = `CIPHERTEXT_WIDTH'd11516263;
cipher_text[122] = `CIPHERTEXT_WIDTH'd11129259;
cipher_text[123] = `CIPHERTEXT_WIDTH'd10446326;
cipher_text[124] = `CIPHERTEXT_WIDTH'd10030738;
cipher_text[125] = `CIPHERTEXT_WIDTH'd12827692;
cipher_text[126] = `CIPHERTEXT_WIDTH'd11282280;
cipher_text[127] = `CIPHERTEXT_WIDTH'd4766930;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 17;
cipher_text[0] = `CIPHERTEXT_WIDTH'd11038724;
cipher_text[1] = `CIPHERTEXT_WIDTH'd4066462;
cipher_text[2] = `CIPHERTEXT_WIDTH'd3253029;
cipher_text[3] = `CIPHERTEXT_WIDTH'd6841616;
cipher_text[4] = `CIPHERTEXT_WIDTH'd5470517;
cipher_text[5] = `CIPHERTEXT_WIDTH'd7037324;
cipher_text[6] = `CIPHERTEXT_WIDTH'd5118189;
cipher_text[7] = `CIPHERTEXT_WIDTH'd8202419;
cipher_text[8] = `CIPHERTEXT_WIDTH'd4562005;
cipher_text[9] = `CIPHERTEXT_WIDTH'd10063419;
cipher_text[10] = `CIPHERTEXT_WIDTH'd115374;
cipher_text[11] = `CIPHERTEXT_WIDTH'd7765238;
cipher_text[12] = `CIPHERTEXT_WIDTH'd9250845;
cipher_text[13] = `CIPHERTEXT_WIDTH'd2060143;
cipher_text[14] = `CIPHERTEXT_WIDTH'd5826816;
cipher_text[15] = `CIPHERTEXT_WIDTH'd15500635;
cipher_text[16] = `CIPHERTEXT_WIDTH'd5649501;
cipher_text[17] = `CIPHERTEXT_WIDTH'd7663853;
cipher_text[18] = `CIPHERTEXT_WIDTH'd13107365;
cipher_text[19] = `CIPHERTEXT_WIDTH'd6500006;
cipher_text[20] = `CIPHERTEXT_WIDTH'd15853046;
cipher_text[21] = `CIPHERTEXT_WIDTH'd4828314;
cipher_text[22] = `CIPHERTEXT_WIDTH'd4444586;
cipher_text[23] = `CIPHERTEXT_WIDTH'd7982356;
cipher_text[24] = `CIPHERTEXT_WIDTH'd13687257;
cipher_text[25] = `CIPHERTEXT_WIDTH'd9395585;
cipher_text[26] = `CIPHERTEXT_WIDTH'd696975;
cipher_text[27] = `CIPHERTEXT_WIDTH'd8165556;
cipher_text[28] = `CIPHERTEXT_WIDTH'd8839233;
cipher_text[29] = `CIPHERTEXT_WIDTH'd11111871;
cipher_text[30] = `CIPHERTEXT_WIDTH'd2312528;
cipher_text[31] = `CIPHERTEXT_WIDTH'd2167717;
cipher_text[32] = `CIPHERTEXT_WIDTH'd5806780;
cipher_text[33] = `CIPHERTEXT_WIDTH'd3449920;
cipher_text[34] = `CIPHERTEXT_WIDTH'd10923517;
cipher_text[35] = `CIPHERTEXT_WIDTH'd10147568;
cipher_text[36] = `CIPHERTEXT_WIDTH'd12472904;
cipher_text[37] = `CIPHERTEXT_WIDTH'd2187977;
cipher_text[38] = `CIPHERTEXT_WIDTH'd13844564;
cipher_text[39] = `CIPHERTEXT_WIDTH'd1030745;
cipher_text[40] = `CIPHERTEXT_WIDTH'd13842500;
cipher_text[41] = `CIPHERTEXT_WIDTH'd2778205;
cipher_text[42] = `CIPHERTEXT_WIDTH'd1450701;
cipher_text[43] = `CIPHERTEXT_WIDTH'd13218778;
cipher_text[44] = `CIPHERTEXT_WIDTH'd2926784;
cipher_text[45] = `CIPHERTEXT_WIDTH'd8511532;
cipher_text[46] = `CIPHERTEXT_WIDTH'd3400858;
cipher_text[47] = `CIPHERTEXT_WIDTH'd3810574;
cipher_text[48] = `CIPHERTEXT_WIDTH'd14859776;
cipher_text[49] = `CIPHERTEXT_WIDTH'd14343721;
cipher_text[50] = `CIPHERTEXT_WIDTH'd1397215;
cipher_text[51] = `CIPHERTEXT_WIDTH'd12645351;
cipher_text[52] = `CIPHERTEXT_WIDTH'd1015492;
cipher_text[53] = `CIPHERTEXT_WIDTH'd7617203;
cipher_text[54] = `CIPHERTEXT_WIDTH'd8663056;
cipher_text[55] = `CIPHERTEXT_WIDTH'd4621068;
cipher_text[56] = `CIPHERTEXT_WIDTH'd13346593;
cipher_text[57] = `CIPHERTEXT_WIDTH'd2502555;
cipher_text[58] = `CIPHERTEXT_WIDTH'd13545134;
cipher_text[59] = `CIPHERTEXT_WIDTH'd7490448;
cipher_text[60] = `CIPHERTEXT_WIDTH'd10052863;
cipher_text[61] = `CIPHERTEXT_WIDTH'd3731001;
cipher_text[62] = `CIPHERTEXT_WIDTH'd16764625;
cipher_text[63] = `CIPHERTEXT_WIDTH'd1715460;
cipher_text[64] = `CIPHERTEXT_WIDTH'd14681085;
cipher_text[65] = `CIPHERTEXT_WIDTH'd7776175;
cipher_text[66] = `CIPHERTEXT_WIDTH'd7117231;
cipher_text[67] = `CIPHERTEXT_WIDTH'd6343682;
cipher_text[68] = `CIPHERTEXT_WIDTH'd8807104;
cipher_text[69] = `CIPHERTEXT_WIDTH'd9319026;
cipher_text[70] = `CIPHERTEXT_WIDTH'd5758013;
cipher_text[71] = `CIPHERTEXT_WIDTH'd3013617;
cipher_text[72] = `CIPHERTEXT_WIDTH'd3393485;
cipher_text[73] = `CIPHERTEXT_WIDTH'd14200308;
cipher_text[74] = `CIPHERTEXT_WIDTH'd10552866;
cipher_text[75] = `CIPHERTEXT_WIDTH'd6548953;
cipher_text[76] = `CIPHERTEXT_WIDTH'd944355;
cipher_text[77] = `CIPHERTEXT_WIDTH'd149747;
cipher_text[78] = `CIPHERTEXT_WIDTH'd12639708;
cipher_text[79] = `CIPHERTEXT_WIDTH'd1760225;
cipher_text[80] = `CIPHERTEXT_WIDTH'd14232382;
cipher_text[81] = `CIPHERTEXT_WIDTH'd15378443;
cipher_text[82] = `CIPHERTEXT_WIDTH'd4871602;
cipher_text[83] = `CIPHERTEXT_WIDTH'd11540423;
cipher_text[84] = `CIPHERTEXT_WIDTH'd4753303;
cipher_text[85] = `CIPHERTEXT_WIDTH'd8039446;
cipher_text[86] = `CIPHERTEXT_WIDTH'd11113076;
cipher_text[87] = `CIPHERTEXT_WIDTH'd11954308;
cipher_text[88] = `CIPHERTEXT_WIDTH'd16716084;
cipher_text[89] = `CIPHERTEXT_WIDTH'd11711608;
cipher_text[90] = `CIPHERTEXT_WIDTH'd1318304;
cipher_text[91] = `CIPHERTEXT_WIDTH'd1982107;
cipher_text[92] = `CIPHERTEXT_WIDTH'd1234933;
cipher_text[93] = `CIPHERTEXT_WIDTH'd14641542;
cipher_text[94] = `CIPHERTEXT_WIDTH'd10055158;
cipher_text[95] = `CIPHERTEXT_WIDTH'd16081224;
cipher_text[96] = `CIPHERTEXT_WIDTH'd5458827;
cipher_text[97] = `CIPHERTEXT_WIDTH'd10223349;
cipher_text[98] = `CIPHERTEXT_WIDTH'd8149105;
cipher_text[99] = `CIPHERTEXT_WIDTH'd9441966;
cipher_text[100] = `CIPHERTEXT_WIDTH'd4286957;
cipher_text[101] = `CIPHERTEXT_WIDTH'd10106250;
cipher_text[102] = `CIPHERTEXT_WIDTH'd7955696;
cipher_text[103] = `CIPHERTEXT_WIDTH'd12516757;
cipher_text[104] = `CIPHERTEXT_WIDTH'd15125796;
cipher_text[105] = `CIPHERTEXT_WIDTH'd1812495;
cipher_text[106] = `CIPHERTEXT_WIDTH'd6692064;
cipher_text[107] = `CIPHERTEXT_WIDTH'd7046809;
cipher_text[108] = `CIPHERTEXT_WIDTH'd4333170;
cipher_text[109] = `CIPHERTEXT_WIDTH'd12479719;
cipher_text[110] = `CIPHERTEXT_WIDTH'd14592059;
cipher_text[111] = `CIPHERTEXT_WIDTH'd2192978;
cipher_text[112] = `CIPHERTEXT_WIDTH'd8209297;
cipher_text[113] = `CIPHERTEXT_WIDTH'd15183386;
cipher_text[114] = `CIPHERTEXT_WIDTH'd15445225;
cipher_text[115] = `CIPHERTEXT_WIDTH'd13313210;
cipher_text[116] = `CIPHERTEXT_WIDTH'd3974768;
cipher_text[117] = `CIPHERTEXT_WIDTH'd9229822;
cipher_text[118] = `CIPHERTEXT_WIDTH'd10052311;
cipher_text[119] = `CIPHERTEXT_WIDTH'd13170379;
cipher_text[120] = `CIPHERTEXT_WIDTH'd2374581;
cipher_text[121] = `CIPHERTEXT_WIDTH'd16045218;
cipher_text[122] = `CIPHERTEXT_WIDTH'd3209590;
cipher_text[123] = `CIPHERTEXT_WIDTH'd3436397;
cipher_text[124] = `CIPHERTEXT_WIDTH'd15931794;
cipher_text[125] = `CIPHERTEXT_WIDTH'd15460152;
cipher_text[126] = `CIPHERTEXT_WIDTH'd7282196;
cipher_text[127] = `CIPHERTEXT_WIDTH'd2750042;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 18;
cipher_text[0] = `CIPHERTEXT_WIDTH'd928541;
cipher_text[1] = `CIPHERTEXT_WIDTH'd8269887;
cipher_text[2] = `CIPHERTEXT_WIDTH'd2357390;
cipher_text[3] = `CIPHERTEXT_WIDTH'd15306697;
cipher_text[4] = `CIPHERTEXT_WIDTH'd14867034;
cipher_text[5] = `CIPHERTEXT_WIDTH'd6755991;
cipher_text[6] = `CIPHERTEXT_WIDTH'd4162141;
cipher_text[7] = `CIPHERTEXT_WIDTH'd5237769;
cipher_text[8] = `CIPHERTEXT_WIDTH'd10820098;
cipher_text[9] = `CIPHERTEXT_WIDTH'd3697026;
cipher_text[10] = `CIPHERTEXT_WIDTH'd3491737;
cipher_text[11] = `CIPHERTEXT_WIDTH'd5739394;
cipher_text[12] = `CIPHERTEXT_WIDTH'd3451461;
cipher_text[13] = `CIPHERTEXT_WIDTH'd2322121;
cipher_text[14] = `CIPHERTEXT_WIDTH'd8978171;
cipher_text[15] = `CIPHERTEXT_WIDTH'd1390473;
cipher_text[16] = `CIPHERTEXT_WIDTH'd4710474;
cipher_text[17] = `CIPHERTEXT_WIDTH'd6617523;
cipher_text[18] = `CIPHERTEXT_WIDTH'd10992776;
cipher_text[19] = `CIPHERTEXT_WIDTH'd16389363;
cipher_text[20] = `CIPHERTEXT_WIDTH'd10433783;
cipher_text[21] = `CIPHERTEXT_WIDTH'd6813223;
cipher_text[22] = `CIPHERTEXT_WIDTH'd16391268;
cipher_text[23] = `CIPHERTEXT_WIDTH'd11718583;
cipher_text[24] = `CIPHERTEXT_WIDTH'd5406859;
cipher_text[25] = `CIPHERTEXT_WIDTH'd8465148;
cipher_text[26] = `CIPHERTEXT_WIDTH'd2131269;
cipher_text[27] = `CIPHERTEXT_WIDTH'd4965471;
cipher_text[28] = `CIPHERTEXT_WIDTH'd7174665;
cipher_text[29] = `CIPHERTEXT_WIDTH'd4222601;
cipher_text[30] = `CIPHERTEXT_WIDTH'd15647755;
cipher_text[31] = `CIPHERTEXT_WIDTH'd701475;
cipher_text[32] = `CIPHERTEXT_WIDTH'd12780423;
cipher_text[33] = `CIPHERTEXT_WIDTH'd7248741;
cipher_text[34] = `CIPHERTEXT_WIDTH'd5465809;
cipher_text[35] = `CIPHERTEXT_WIDTH'd6859450;
cipher_text[36] = `CIPHERTEXT_WIDTH'd15160959;
cipher_text[37] = `CIPHERTEXT_WIDTH'd6739888;
cipher_text[38] = `CIPHERTEXT_WIDTH'd4672204;
cipher_text[39] = `CIPHERTEXT_WIDTH'd11074615;
cipher_text[40] = `CIPHERTEXT_WIDTH'd596922;
cipher_text[41] = `CIPHERTEXT_WIDTH'd16208039;
cipher_text[42] = `CIPHERTEXT_WIDTH'd9537804;
cipher_text[43] = `CIPHERTEXT_WIDTH'd13419799;
cipher_text[44] = `CIPHERTEXT_WIDTH'd9336044;
cipher_text[45] = `CIPHERTEXT_WIDTH'd16528003;
cipher_text[46] = `CIPHERTEXT_WIDTH'd5797343;
cipher_text[47] = `CIPHERTEXT_WIDTH'd9932999;
cipher_text[48] = `CIPHERTEXT_WIDTH'd10282782;
cipher_text[49] = `CIPHERTEXT_WIDTH'd12952163;
cipher_text[50] = `CIPHERTEXT_WIDTH'd7998042;
cipher_text[51] = `CIPHERTEXT_WIDTH'd10895739;
cipher_text[52] = `CIPHERTEXT_WIDTH'd5377722;
cipher_text[53] = `CIPHERTEXT_WIDTH'd15971945;
cipher_text[54] = `CIPHERTEXT_WIDTH'd11357769;
cipher_text[55] = `CIPHERTEXT_WIDTH'd4308641;
cipher_text[56] = `CIPHERTEXT_WIDTH'd6104132;
cipher_text[57] = `CIPHERTEXT_WIDTH'd6712380;
cipher_text[58] = `CIPHERTEXT_WIDTH'd10373925;
cipher_text[59] = `CIPHERTEXT_WIDTH'd2705481;
cipher_text[60] = `CIPHERTEXT_WIDTH'd5600920;
cipher_text[61] = `CIPHERTEXT_WIDTH'd7405983;
cipher_text[62] = `CIPHERTEXT_WIDTH'd9637814;
cipher_text[63] = `CIPHERTEXT_WIDTH'd12811505;
cipher_text[64] = `CIPHERTEXT_WIDTH'd11688113;
cipher_text[65] = `CIPHERTEXT_WIDTH'd7803695;
cipher_text[66] = `CIPHERTEXT_WIDTH'd9652337;
cipher_text[67] = `CIPHERTEXT_WIDTH'd312518;
cipher_text[68] = `CIPHERTEXT_WIDTH'd12882468;
cipher_text[69] = `CIPHERTEXT_WIDTH'd7386733;
cipher_text[70] = `CIPHERTEXT_WIDTH'd4457039;
cipher_text[71] = `CIPHERTEXT_WIDTH'd15022146;
cipher_text[72] = `CIPHERTEXT_WIDTH'd2533961;
cipher_text[73] = `CIPHERTEXT_WIDTH'd12928132;
cipher_text[74] = `CIPHERTEXT_WIDTH'd580595;
cipher_text[75] = `CIPHERTEXT_WIDTH'd7665841;
cipher_text[76] = `CIPHERTEXT_WIDTH'd7934233;
cipher_text[77] = `CIPHERTEXT_WIDTH'd13917490;
cipher_text[78] = `CIPHERTEXT_WIDTH'd1141072;
cipher_text[79] = `CIPHERTEXT_WIDTH'd15453003;
cipher_text[80] = `CIPHERTEXT_WIDTH'd11463955;
cipher_text[81] = `CIPHERTEXT_WIDTH'd6818533;
cipher_text[82] = `CIPHERTEXT_WIDTH'd11103208;
cipher_text[83] = `CIPHERTEXT_WIDTH'd15749008;
cipher_text[84] = `CIPHERTEXT_WIDTH'd7302741;
cipher_text[85] = `CIPHERTEXT_WIDTH'd2382387;
cipher_text[86] = `CIPHERTEXT_WIDTH'd12304731;
cipher_text[87] = `CIPHERTEXT_WIDTH'd3217454;
cipher_text[88] = `CIPHERTEXT_WIDTH'd5835063;
cipher_text[89] = `CIPHERTEXT_WIDTH'd6696512;
cipher_text[90] = `CIPHERTEXT_WIDTH'd4450509;
cipher_text[91] = `CIPHERTEXT_WIDTH'd10625840;
cipher_text[92] = `CIPHERTEXT_WIDTH'd8333876;
cipher_text[93] = `CIPHERTEXT_WIDTH'd3922801;
cipher_text[94] = `CIPHERTEXT_WIDTH'd15398353;
cipher_text[95] = `CIPHERTEXT_WIDTH'd14408231;
cipher_text[96] = `CIPHERTEXT_WIDTH'd14432529;
cipher_text[97] = `CIPHERTEXT_WIDTH'd9555359;
cipher_text[98] = `CIPHERTEXT_WIDTH'd8600087;
cipher_text[99] = `CIPHERTEXT_WIDTH'd13826120;
cipher_text[100] = `CIPHERTEXT_WIDTH'd9452549;
cipher_text[101] = `CIPHERTEXT_WIDTH'd13153156;
cipher_text[102] = `CIPHERTEXT_WIDTH'd11152173;
cipher_text[103] = `CIPHERTEXT_WIDTH'd13673233;
cipher_text[104] = `CIPHERTEXT_WIDTH'd10409615;
cipher_text[105] = `CIPHERTEXT_WIDTH'd8783248;
cipher_text[106] = `CIPHERTEXT_WIDTH'd7003437;
cipher_text[107] = `CIPHERTEXT_WIDTH'd15133459;
cipher_text[108] = `CIPHERTEXT_WIDTH'd5739309;
cipher_text[109] = `CIPHERTEXT_WIDTH'd5887391;
cipher_text[110] = `CIPHERTEXT_WIDTH'd7022904;
cipher_text[111] = `CIPHERTEXT_WIDTH'd3537368;
cipher_text[112] = `CIPHERTEXT_WIDTH'd3863149;
cipher_text[113] = `CIPHERTEXT_WIDTH'd14330480;
cipher_text[114] = `CIPHERTEXT_WIDTH'd10416237;
cipher_text[115] = `CIPHERTEXT_WIDTH'd2895472;
cipher_text[116] = `CIPHERTEXT_WIDTH'd9125571;
cipher_text[117] = `CIPHERTEXT_WIDTH'd16003504;
cipher_text[118] = `CIPHERTEXT_WIDTH'd7779555;
cipher_text[119] = `CIPHERTEXT_WIDTH'd11876425;
cipher_text[120] = `CIPHERTEXT_WIDTH'd6311452;
cipher_text[121] = `CIPHERTEXT_WIDTH'd5178889;
cipher_text[122] = `CIPHERTEXT_WIDTH'd12885706;
cipher_text[123] = `CIPHERTEXT_WIDTH'd599916;
cipher_text[124] = `CIPHERTEXT_WIDTH'd1425569;
cipher_text[125] = `CIPHERTEXT_WIDTH'd14875817;
cipher_text[126] = `CIPHERTEXT_WIDTH'd1899563;
cipher_text[127] = `CIPHERTEXT_WIDTH'd15348220;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 19;
cipher_text[0] = `CIPHERTEXT_WIDTH'd14185663;
cipher_text[1] = `CIPHERTEXT_WIDTH'd5663038;
cipher_text[2] = `CIPHERTEXT_WIDTH'd11968153;
cipher_text[3] = `CIPHERTEXT_WIDTH'd13796964;
cipher_text[4] = `CIPHERTEXT_WIDTH'd1049579;
cipher_text[5] = `CIPHERTEXT_WIDTH'd2463395;
cipher_text[6] = `CIPHERTEXT_WIDTH'd12731406;
cipher_text[7] = `CIPHERTEXT_WIDTH'd4044761;
cipher_text[8] = `CIPHERTEXT_WIDTH'd15067765;
cipher_text[9] = `CIPHERTEXT_WIDTH'd13435001;
cipher_text[10] = `CIPHERTEXT_WIDTH'd9547042;
cipher_text[11] = `CIPHERTEXT_WIDTH'd7377775;
cipher_text[12] = `CIPHERTEXT_WIDTH'd11093818;
cipher_text[13] = `CIPHERTEXT_WIDTH'd5095149;
cipher_text[14] = `CIPHERTEXT_WIDTH'd9807085;
cipher_text[15] = `CIPHERTEXT_WIDTH'd14690010;
cipher_text[16] = `CIPHERTEXT_WIDTH'd2996333;
cipher_text[17] = `CIPHERTEXT_WIDTH'd4579896;
cipher_text[18] = `CIPHERTEXT_WIDTH'd6879527;
cipher_text[19] = `CIPHERTEXT_WIDTH'd498529;
cipher_text[20] = `CIPHERTEXT_WIDTH'd9834814;
cipher_text[21] = `CIPHERTEXT_WIDTH'd7945603;
cipher_text[22] = `CIPHERTEXT_WIDTH'd6581970;
cipher_text[23] = `CIPHERTEXT_WIDTH'd8218935;
cipher_text[24] = `CIPHERTEXT_WIDTH'd5359670;
cipher_text[25] = `CIPHERTEXT_WIDTH'd10214005;
cipher_text[26] = `CIPHERTEXT_WIDTH'd7700427;
cipher_text[27] = `CIPHERTEXT_WIDTH'd10579263;
cipher_text[28] = `CIPHERTEXT_WIDTH'd1644355;
cipher_text[29] = `CIPHERTEXT_WIDTH'd14586619;
cipher_text[30] = `CIPHERTEXT_WIDTH'd7052437;
cipher_text[31] = `CIPHERTEXT_WIDTH'd13296967;
cipher_text[32] = `CIPHERTEXT_WIDTH'd6726898;
cipher_text[33] = `CIPHERTEXT_WIDTH'd14841350;
cipher_text[34] = `CIPHERTEXT_WIDTH'd16545527;
cipher_text[35] = `CIPHERTEXT_WIDTH'd13605601;
cipher_text[36] = `CIPHERTEXT_WIDTH'd6516064;
cipher_text[37] = `CIPHERTEXT_WIDTH'd9157904;
cipher_text[38] = `CIPHERTEXT_WIDTH'd13418233;
cipher_text[39] = `CIPHERTEXT_WIDTH'd6701913;
cipher_text[40] = `CIPHERTEXT_WIDTH'd15160282;
cipher_text[41] = `CIPHERTEXT_WIDTH'd8807803;
cipher_text[42] = `CIPHERTEXT_WIDTH'd5674680;
cipher_text[43] = `CIPHERTEXT_WIDTH'd3184366;
cipher_text[44] = `CIPHERTEXT_WIDTH'd1204734;
cipher_text[45] = `CIPHERTEXT_WIDTH'd9771692;
cipher_text[46] = `CIPHERTEXT_WIDTH'd3794881;
cipher_text[47] = `CIPHERTEXT_WIDTH'd4881584;
cipher_text[48] = `CIPHERTEXT_WIDTH'd7354217;
cipher_text[49] = `CIPHERTEXT_WIDTH'd7922569;
cipher_text[50] = `CIPHERTEXT_WIDTH'd16281576;
cipher_text[51] = `CIPHERTEXT_WIDTH'd2231625;
cipher_text[52] = `CIPHERTEXT_WIDTH'd16525950;
cipher_text[53] = `CIPHERTEXT_WIDTH'd11445675;
cipher_text[54] = `CIPHERTEXT_WIDTH'd3355899;
cipher_text[55] = `CIPHERTEXT_WIDTH'd14166200;
cipher_text[56] = `CIPHERTEXT_WIDTH'd2394602;
cipher_text[57] = `CIPHERTEXT_WIDTH'd13095394;
cipher_text[58] = `CIPHERTEXT_WIDTH'd7798602;
cipher_text[59] = `CIPHERTEXT_WIDTH'd3188248;
cipher_text[60] = `CIPHERTEXT_WIDTH'd16605162;
cipher_text[61] = `CIPHERTEXT_WIDTH'd11972825;
cipher_text[62] = `CIPHERTEXT_WIDTH'd15968155;
cipher_text[63] = `CIPHERTEXT_WIDTH'd1213052;
cipher_text[64] = `CIPHERTEXT_WIDTH'd12167754;
cipher_text[65] = `CIPHERTEXT_WIDTH'd15294891;
cipher_text[66] = `CIPHERTEXT_WIDTH'd1023272;
cipher_text[67] = `CIPHERTEXT_WIDTH'd9164270;
cipher_text[68] = `CIPHERTEXT_WIDTH'd15124425;
cipher_text[69] = `CIPHERTEXT_WIDTH'd7795621;
cipher_text[70] = `CIPHERTEXT_WIDTH'd6879609;
cipher_text[71] = `CIPHERTEXT_WIDTH'd6725035;
cipher_text[72] = `CIPHERTEXT_WIDTH'd13099823;
cipher_text[73] = `CIPHERTEXT_WIDTH'd1688074;
cipher_text[74] = `CIPHERTEXT_WIDTH'd3167734;
cipher_text[75] = `CIPHERTEXT_WIDTH'd16271167;
cipher_text[76] = `CIPHERTEXT_WIDTH'd10059979;
cipher_text[77] = `CIPHERTEXT_WIDTH'd5191247;
cipher_text[78] = `CIPHERTEXT_WIDTH'd10611919;
cipher_text[79] = `CIPHERTEXT_WIDTH'd9967758;
cipher_text[80] = `CIPHERTEXT_WIDTH'd11450704;
cipher_text[81] = `CIPHERTEXT_WIDTH'd7144729;
cipher_text[82] = `CIPHERTEXT_WIDTH'd5398147;
cipher_text[83] = `CIPHERTEXT_WIDTH'd7973302;
cipher_text[84] = `CIPHERTEXT_WIDTH'd15917019;
cipher_text[85] = `CIPHERTEXT_WIDTH'd3764938;
cipher_text[86] = `CIPHERTEXT_WIDTH'd7628434;
cipher_text[87] = `CIPHERTEXT_WIDTH'd3127191;
cipher_text[88] = `CIPHERTEXT_WIDTH'd15905739;
cipher_text[89] = `CIPHERTEXT_WIDTH'd15982318;
cipher_text[90] = `CIPHERTEXT_WIDTH'd12150372;
cipher_text[91] = `CIPHERTEXT_WIDTH'd11251850;
cipher_text[92] = `CIPHERTEXT_WIDTH'd3877509;
cipher_text[93] = `CIPHERTEXT_WIDTH'd11234292;
cipher_text[94] = `CIPHERTEXT_WIDTH'd2352101;
cipher_text[95] = `CIPHERTEXT_WIDTH'd1535545;
cipher_text[96] = `CIPHERTEXT_WIDTH'd3144823;
cipher_text[97] = `CIPHERTEXT_WIDTH'd9170918;
cipher_text[98] = `CIPHERTEXT_WIDTH'd10259182;
cipher_text[99] = `CIPHERTEXT_WIDTH'd16473610;
cipher_text[100] = `CIPHERTEXT_WIDTH'd2444509;
cipher_text[101] = `CIPHERTEXT_WIDTH'd10842899;
cipher_text[102] = `CIPHERTEXT_WIDTH'd10117191;
cipher_text[103] = `CIPHERTEXT_WIDTH'd1185292;
cipher_text[104] = `CIPHERTEXT_WIDTH'd558475;
cipher_text[105] = `CIPHERTEXT_WIDTH'd4854333;
cipher_text[106] = `CIPHERTEXT_WIDTH'd11871624;
cipher_text[107] = `CIPHERTEXT_WIDTH'd3809158;
cipher_text[108] = `CIPHERTEXT_WIDTH'd5775671;
cipher_text[109] = `CIPHERTEXT_WIDTH'd13113567;
cipher_text[110] = `CIPHERTEXT_WIDTH'd4375580;
cipher_text[111] = `CIPHERTEXT_WIDTH'd3660658;
cipher_text[112] = `CIPHERTEXT_WIDTH'd9104505;
cipher_text[113] = `CIPHERTEXT_WIDTH'd8144247;
cipher_text[114] = `CIPHERTEXT_WIDTH'd8822254;
cipher_text[115] = `CIPHERTEXT_WIDTH'd11488438;
cipher_text[116] = `CIPHERTEXT_WIDTH'd10713074;
cipher_text[117] = `CIPHERTEXT_WIDTH'd13995724;
cipher_text[118] = `CIPHERTEXT_WIDTH'd10047561;
cipher_text[119] = `CIPHERTEXT_WIDTH'd10625191;
cipher_text[120] = `CIPHERTEXT_WIDTH'd16292271;
cipher_text[121] = `CIPHERTEXT_WIDTH'd834371;
cipher_text[122] = `CIPHERTEXT_WIDTH'd6920466;
cipher_text[123] = `CIPHERTEXT_WIDTH'd4381345;
cipher_text[124] = `CIPHERTEXT_WIDTH'd16021488;
cipher_text[125] = `CIPHERTEXT_WIDTH'd13253297;
cipher_text[126] = `CIPHERTEXT_WIDTH'd7712061;
cipher_text[127] = `CIPHERTEXT_WIDTH'd10496012;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 20;
cipher_text[0] = `CIPHERTEXT_WIDTH'd16728946;
cipher_text[1] = `CIPHERTEXT_WIDTH'd15342517;
cipher_text[2] = `CIPHERTEXT_WIDTH'd3526956;
cipher_text[3] = `CIPHERTEXT_WIDTH'd11597309;
cipher_text[4] = `CIPHERTEXT_WIDTH'd9357569;
cipher_text[5] = `CIPHERTEXT_WIDTH'd3729319;
cipher_text[6] = `CIPHERTEXT_WIDTH'd16601350;
cipher_text[7] = `CIPHERTEXT_WIDTH'd15372332;
cipher_text[8] = `CIPHERTEXT_WIDTH'd6650452;
cipher_text[9] = `CIPHERTEXT_WIDTH'd15036065;
cipher_text[10] = `CIPHERTEXT_WIDTH'd3232867;
cipher_text[11] = `CIPHERTEXT_WIDTH'd7955396;
cipher_text[12] = `CIPHERTEXT_WIDTH'd11365371;
cipher_text[13] = `CIPHERTEXT_WIDTH'd5106508;
cipher_text[14] = `CIPHERTEXT_WIDTH'd13602347;
cipher_text[15] = `CIPHERTEXT_WIDTH'd13452847;
cipher_text[16] = `CIPHERTEXT_WIDTH'd1991814;
cipher_text[17] = `CIPHERTEXT_WIDTH'd3070531;
cipher_text[18] = `CIPHERTEXT_WIDTH'd12554274;
cipher_text[19] = `CIPHERTEXT_WIDTH'd11114235;
cipher_text[20] = `CIPHERTEXT_WIDTH'd15668113;
cipher_text[21] = `CIPHERTEXT_WIDTH'd13333782;
cipher_text[22] = `CIPHERTEXT_WIDTH'd9635116;
cipher_text[23] = `CIPHERTEXT_WIDTH'd1476233;
cipher_text[24] = `CIPHERTEXT_WIDTH'd10268759;
cipher_text[25] = `CIPHERTEXT_WIDTH'd10571594;
cipher_text[26] = `CIPHERTEXT_WIDTH'd15323998;
cipher_text[27] = `CIPHERTEXT_WIDTH'd4522239;
cipher_text[28] = `CIPHERTEXT_WIDTH'd16522097;
cipher_text[29] = `CIPHERTEXT_WIDTH'd13408722;
cipher_text[30] = `CIPHERTEXT_WIDTH'd4168060;
cipher_text[31] = `CIPHERTEXT_WIDTH'd5209844;
cipher_text[32] = `CIPHERTEXT_WIDTH'd149887;
cipher_text[33] = `CIPHERTEXT_WIDTH'd1886930;
cipher_text[34] = `CIPHERTEXT_WIDTH'd6475351;
cipher_text[35] = `CIPHERTEXT_WIDTH'd15248632;
cipher_text[36] = `CIPHERTEXT_WIDTH'd13798942;
cipher_text[37] = `CIPHERTEXT_WIDTH'd3473633;
cipher_text[38] = `CIPHERTEXT_WIDTH'd6974523;
cipher_text[39] = `CIPHERTEXT_WIDTH'd9376546;
cipher_text[40] = `CIPHERTEXT_WIDTH'd12376840;
cipher_text[41] = `CIPHERTEXT_WIDTH'd5287989;
cipher_text[42] = `CIPHERTEXT_WIDTH'd11710105;
cipher_text[43] = `CIPHERTEXT_WIDTH'd11783612;
cipher_text[44] = `CIPHERTEXT_WIDTH'd15750236;
cipher_text[45] = `CIPHERTEXT_WIDTH'd16647015;
cipher_text[46] = `CIPHERTEXT_WIDTH'd3671119;
cipher_text[47] = `CIPHERTEXT_WIDTH'd10396478;
cipher_text[48] = `CIPHERTEXT_WIDTH'd772631;
cipher_text[49] = `CIPHERTEXT_WIDTH'd5843538;
cipher_text[50] = `CIPHERTEXT_WIDTH'd1328990;
cipher_text[51] = `CIPHERTEXT_WIDTH'd4404588;
cipher_text[52] = `CIPHERTEXT_WIDTH'd15758404;
cipher_text[53] = `CIPHERTEXT_WIDTH'd14746588;
cipher_text[54] = `CIPHERTEXT_WIDTH'd2472683;
cipher_text[55] = `CIPHERTEXT_WIDTH'd2681406;
cipher_text[56] = `CIPHERTEXT_WIDTH'd7698548;
cipher_text[57] = `CIPHERTEXT_WIDTH'd14626768;
cipher_text[58] = `CIPHERTEXT_WIDTH'd1382509;
cipher_text[59] = `CIPHERTEXT_WIDTH'd1135275;
cipher_text[60] = `CIPHERTEXT_WIDTH'd15304777;
cipher_text[61] = `CIPHERTEXT_WIDTH'd10446061;
cipher_text[62] = `CIPHERTEXT_WIDTH'd13891912;
cipher_text[63] = `CIPHERTEXT_WIDTH'd5899497;
cipher_text[64] = `CIPHERTEXT_WIDTH'd5420540;
cipher_text[65] = `CIPHERTEXT_WIDTH'd1515213;
cipher_text[66] = `CIPHERTEXT_WIDTH'd2636896;
cipher_text[67] = `CIPHERTEXT_WIDTH'd9260013;
cipher_text[68] = `CIPHERTEXT_WIDTH'd15099056;
cipher_text[69] = `CIPHERTEXT_WIDTH'd6823973;
cipher_text[70] = `CIPHERTEXT_WIDTH'd11180510;
cipher_text[71] = `CIPHERTEXT_WIDTH'd6749925;
cipher_text[72] = `CIPHERTEXT_WIDTH'd11618616;
cipher_text[73] = `CIPHERTEXT_WIDTH'd12647034;
cipher_text[74] = `CIPHERTEXT_WIDTH'd4536440;
cipher_text[75] = `CIPHERTEXT_WIDTH'd2102545;
cipher_text[76] = `CIPHERTEXT_WIDTH'd3444425;
cipher_text[77] = `CIPHERTEXT_WIDTH'd15005274;
cipher_text[78] = `CIPHERTEXT_WIDTH'd11594000;
cipher_text[79] = `CIPHERTEXT_WIDTH'd8141444;
cipher_text[80] = `CIPHERTEXT_WIDTH'd9866533;
cipher_text[81] = `CIPHERTEXT_WIDTH'd16355097;
cipher_text[82] = `CIPHERTEXT_WIDTH'd14681001;
cipher_text[83] = `CIPHERTEXT_WIDTH'd304717;
cipher_text[84] = `CIPHERTEXT_WIDTH'd16351333;
cipher_text[85] = `CIPHERTEXT_WIDTH'd8371349;
cipher_text[86] = `CIPHERTEXT_WIDTH'd16560107;
cipher_text[87] = `CIPHERTEXT_WIDTH'd6329614;
cipher_text[88] = `CIPHERTEXT_WIDTH'd10142569;
cipher_text[89] = `CIPHERTEXT_WIDTH'd5636754;
cipher_text[90] = `CIPHERTEXT_WIDTH'd11781435;
cipher_text[91] = `CIPHERTEXT_WIDTH'd1180453;
cipher_text[92] = `CIPHERTEXT_WIDTH'd10299499;
cipher_text[93] = `CIPHERTEXT_WIDTH'd2453942;
cipher_text[94] = `CIPHERTEXT_WIDTH'd6515789;
cipher_text[95] = `CIPHERTEXT_WIDTH'd12678354;
cipher_text[96] = `CIPHERTEXT_WIDTH'd13415917;
cipher_text[97] = `CIPHERTEXT_WIDTH'd7077797;
cipher_text[98] = `CIPHERTEXT_WIDTH'd5093630;
cipher_text[99] = `CIPHERTEXT_WIDTH'd12407857;
cipher_text[100] = `CIPHERTEXT_WIDTH'd6131084;
cipher_text[101] = `CIPHERTEXT_WIDTH'd2888822;
cipher_text[102] = `CIPHERTEXT_WIDTH'd4623947;
cipher_text[103] = `CIPHERTEXT_WIDTH'd15917737;
cipher_text[104] = `CIPHERTEXT_WIDTH'd4899113;
cipher_text[105] = `CIPHERTEXT_WIDTH'd11207442;
cipher_text[106] = `CIPHERTEXT_WIDTH'd1308047;
cipher_text[107] = `CIPHERTEXT_WIDTH'd2947530;
cipher_text[108] = `CIPHERTEXT_WIDTH'd10903467;
cipher_text[109] = `CIPHERTEXT_WIDTH'd11629952;
cipher_text[110] = `CIPHERTEXT_WIDTH'd5830762;
cipher_text[111] = `CIPHERTEXT_WIDTH'd13387825;
cipher_text[112] = `CIPHERTEXT_WIDTH'd8702680;
cipher_text[113] = `CIPHERTEXT_WIDTH'd10975965;
cipher_text[114] = `CIPHERTEXT_WIDTH'd12880413;
cipher_text[115] = `CIPHERTEXT_WIDTH'd11121843;
cipher_text[116] = `CIPHERTEXT_WIDTH'd3064667;
cipher_text[117] = `CIPHERTEXT_WIDTH'd14861075;
cipher_text[118] = `CIPHERTEXT_WIDTH'd3567089;
cipher_text[119] = `CIPHERTEXT_WIDTH'd16575206;
cipher_text[120] = `CIPHERTEXT_WIDTH'd9469529;
cipher_text[121] = `CIPHERTEXT_WIDTH'd9543193;
cipher_text[122] = `CIPHERTEXT_WIDTH'd11072024;
cipher_text[123] = `CIPHERTEXT_WIDTH'd11980178;
cipher_text[124] = `CIPHERTEXT_WIDTH'd12621677;
cipher_text[125] = `CIPHERTEXT_WIDTH'd4981026;
cipher_text[126] = `CIPHERTEXT_WIDTH'd14133940;
cipher_text[127] = `CIPHERTEXT_WIDTH'd1880284;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 21;
cipher_text[0] = `CIPHERTEXT_WIDTH'd7478705;
cipher_text[1] = `CIPHERTEXT_WIDTH'd2809753;
cipher_text[2] = `CIPHERTEXT_WIDTH'd5962396;
cipher_text[3] = `CIPHERTEXT_WIDTH'd3695357;
cipher_text[4] = `CIPHERTEXT_WIDTH'd16570663;
cipher_text[5] = `CIPHERTEXT_WIDTH'd7324647;
cipher_text[6] = `CIPHERTEXT_WIDTH'd10472732;
cipher_text[7] = `CIPHERTEXT_WIDTH'd1009914;
cipher_text[8] = `CIPHERTEXT_WIDTH'd6076545;
cipher_text[9] = `CIPHERTEXT_WIDTH'd5154116;
cipher_text[10] = `CIPHERTEXT_WIDTH'd6875867;
cipher_text[11] = `CIPHERTEXT_WIDTH'd9650698;
cipher_text[12] = `CIPHERTEXT_WIDTH'd6123983;
cipher_text[13] = `CIPHERTEXT_WIDTH'd12639373;
cipher_text[14] = `CIPHERTEXT_WIDTH'd1458058;
cipher_text[15] = `CIPHERTEXT_WIDTH'd4543088;
cipher_text[16] = `CIPHERTEXT_WIDTH'd10492233;
cipher_text[17] = `CIPHERTEXT_WIDTH'd8815187;
cipher_text[18] = `CIPHERTEXT_WIDTH'd14659013;
cipher_text[19] = `CIPHERTEXT_WIDTH'd9087487;
cipher_text[20] = `CIPHERTEXT_WIDTH'd10351329;
cipher_text[21] = `CIPHERTEXT_WIDTH'd10364077;
cipher_text[22] = `CIPHERTEXT_WIDTH'd2243953;
cipher_text[23] = `CIPHERTEXT_WIDTH'd3965287;
cipher_text[24] = `CIPHERTEXT_WIDTH'd6773652;
cipher_text[25] = `CIPHERTEXT_WIDTH'd4579442;
cipher_text[26] = `CIPHERTEXT_WIDTH'd3696076;
cipher_text[27] = `CIPHERTEXT_WIDTH'd7889184;
cipher_text[28] = `CIPHERTEXT_WIDTH'd11522819;
cipher_text[29] = `CIPHERTEXT_WIDTH'd12921037;
cipher_text[30] = `CIPHERTEXT_WIDTH'd12611599;
cipher_text[31] = `CIPHERTEXT_WIDTH'd5441881;
cipher_text[32] = `CIPHERTEXT_WIDTH'd9135640;
cipher_text[33] = `CIPHERTEXT_WIDTH'd3440063;
cipher_text[34] = `CIPHERTEXT_WIDTH'd11827105;
cipher_text[35] = `CIPHERTEXT_WIDTH'd7873024;
cipher_text[36] = `CIPHERTEXT_WIDTH'd2515299;
cipher_text[37] = `CIPHERTEXT_WIDTH'd4726834;
cipher_text[38] = `CIPHERTEXT_WIDTH'd7561810;
cipher_text[39] = `CIPHERTEXT_WIDTH'd3332814;
cipher_text[40] = `CIPHERTEXT_WIDTH'd16378900;
cipher_text[41] = `CIPHERTEXT_WIDTH'd8605401;
cipher_text[42] = `CIPHERTEXT_WIDTH'd9106528;
cipher_text[43] = `CIPHERTEXT_WIDTH'd12696340;
cipher_text[44] = `CIPHERTEXT_WIDTH'd6112129;
cipher_text[45] = `CIPHERTEXT_WIDTH'd10535598;
cipher_text[46] = `CIPHERTEXT_WIDTH'd2981584;
cipher_text[47] = `CIPHERTEXT_WIDTH'd6368337;
cipher_text[48] = `CIPHERTEXT_WIDTH'd7587426;
cipher_text[49] = `CIPHERTEXT_WIDTH'd957129;
cipher_text[50] = `CIPHERTEXT_WIDTH'd5449695;
cipher_text[51] = `CIPHERTEXT_WIDTH'd15460442;
cipher_text[52] = `CIPHERTEXT_WIDTH'd1776049;
cipher_text[53] = `CIPHERTEXT_WIDTH'd12970058;
cipher_text[54] = `CIPHERTEXT_WIDTH'd1871682;
cipher_text[55] = `CIPHERTEXT_WIDTH'd8184828;
cipher_text[56] = `CIPHERTEXT_WIDTH'd1685900;
cipher_text[57] = `CIPHERTEXT_WIDTH'd234546;
cipher_text[58] = `CIPHERTEXT_WIDTH'd3355213;
cipher_text[59] = `CIPHERTEXT_WIDTH'd8381046;
cipher_text[60] = `CIPHERTEXT_WIDTH'd8632080;
cipher_text[61] = `CIPHERTEXT_WIDTH'd9723845;
cipher_text[62] = `CIPHERTEXT_WIDTH'd3664116;
cipher_text[63] = `CIPHERTEXT_WIDTH'd12844175;
cipher_text[64] = `CIPHERTEXT_WIDTH'd517921;
cipher_text[65] = `CIPHERTEXT_WIDTH'd8110122;
cipher_text[66] = `CIPHERTEXT_WIDTH'd1033727;
cipher_text[67] = `CIPHERTEXT_WIDTH'd11976307;
cipher_text[68] = `CIPHERTEXT_WIDTH'd15695640;
cipher_text[69] = `CIPHERTEXT_WIDTH'd4366860;
cipher_text[70] = `CIPHERTEXT_WIDTH'd13387714;
cipher_text[71] = `CIPHERTEXT_WIDTH'd9608547;
cipher_text[72] = `CIPHERTEXT_WIDTH'd12721157;
cipher_text[73] = `CIPHERTEXT_WIDTH'd12292029;
cipher_text[74] = `CIPHERTEXT_WIDTH'd4801790;
cipher_text[75] = `CIPHERTEXT_WIDTH'd9326107;
cipher_text[76] = `CIPHERTEXT_WIDTH'd10428758;
cipher_text[77] = `CIPHERTEXT_WIDTH'd9566395;
cipher_text[78] = `CIPHERTEXT_WIDTH'd9801934;
cipher_text[79] = `CIPHERTEXT_WIDTH'd1186425;
cipher_text[80] = `CIPHERTEXT_WIDTH'd3779752;
cipher_text[81] = `CIPHERTEXT_WIDTH'd11638803;
cipher_text[82] = `CIPHERTEXT_WIDTH'd1470446;
cipher_text[83] = `CIPHERTEXT_WIDTH'd13408073;
cipher_text[84] = `CIPHERTEXT_WIDTH'd1980744;
cipher_text[85] = `CIPHERTEXT_WIDTH'd15586188;
cipher_text[86] = `CIPHERTEXT_WIDTH'd11488478;
cipher_text[87] = `CIPHERTEXT_WIDTH'd9454985;
cipher_text[88] = `CIPHERTEXT_WIDTH'd2932991;
cipher_text[89] = `CIPHERTEXT_WIDTH'd9917607;
cipher_text[90] = `CIPHERTEXT_WIDTH'd13877504;
cipher_text[91] = `CIPHERTEXT_WIDTH'd8111967;
cipher_text[92] = `CIPHERTEXT_WIDTH'd13109619;
cipher_text[93] = `CIPHERTEXT_WIDTH'd2395434;
cipher_text[94] = `CIPHERTEXT_WIDTH'd9152666;
cipher_text[95] = `CIPHERTEXT_WIDTH'd11374128;
cipher_text[96] = `CIPHERTEXT_WIDTH'd7865748;
cipher_text[97] = `CIPHERTEXT_WIDTH'd1875527;
cipher_text[98] = `CIPHERTEXT_WIDTH'd9134889;
cipher_text[99] = `CIPHERTEXT_WIDTH'd8977164;
cipher_text[100] = `CIPHERTEXT_WIDTH'd9549273;
cipher_text[101] = `CIPHERTEXT_WIDTH'd15689705;
cipher_text[102] = `CIPHERTEXT_WIDTH'd11701872;
cipher_text[103] = `CIPHERTEXT_WIDTH'd7188111;
cipher_text[104] = `CIPHERTEXT_WIDTH'd15377868;
cipher_text[105] = `CIPHERTEXT_WIDTH'd7585434;
cipher_text[106] = `CIPHERTEXT_WIDTH'd6583135;
cipher_text[107] = `CIPHERTEXT_WIDTH'd5186893;
cipher_text[108] = `CIPHERTEXT_WIDTH'd40567;
cipher_text[109] = `CIPHERTEXT_WIDTH'd6771536;
cipher_text[110] = `CIPHERTEXT_WIDTH'd3999163;
cipher_text[111] = `CIPHERTEXT_WIDTH'd6586821;
cipher_text[112] = `CIPHERTEXT_WIDTH'd14278752;
cipher_text[113] = `CIPHERTEXT_WIDTH'd3851616;
cipher_text[114] = `CIPHERTEXT_WIDTH'd4739660;
cipher_text[115] = `CIPHERTEXT_WIDTH'd8740310;
cipher_text[116] = `CIPHERTEXT_WIDTH'd448431;
cipher_text[117] = `CIPHERTEXT_WIDTH'd7606827;
cipher_text[118] = `CIPHERTEXT_WIDTH'd3433094;
cipher_text[119] = `CIPHERTEXT_WIDTH'd2286612;
cipher_text[120] = `CIPHERTEXT_WIDTH'd7656836;
cipher_text[121] = `CIPHERTEXT_WIDTH'd16296482;
cipher_text[122] = `CIPHERTEXT_WIDTH'd14538777;
cipher_text[123] = `CIPHERTEXT_WIDTH'd1932920;
cipher_text[124] = `CIPHERTEXT_WIDTH'd8552800;
cipher_text[125] = `CIPHERTEXT_WIDTH'd14619019;
cipher_text[126] = `CIPHERTEXT_WIDTH'd4936084;
cipher_text[127] = `CIPHERTEXT_WIDTH'd9193182;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 22;
cipher_text[0] = `CIPHERTEXT_WIDTH'd402377;
cipher_text[1] = `CIPHERTEXT_WIDTH'd15092312;
cipher_text[2] = `CIPHERTEXT_WIDTH'd14402181;
cipher_text[3] = `CIPHERTEXT_WIDTH'd9348985;
cipher_text[4] = `CIPHERTEXT_WIDTH'd13473318;
cipher_text[5] = `CIPHERTEXT_WIDTH'd1497653;
cipher_text[6] = `CIPHERTEXT_WIDTH'd16634400;
cipher_text[7] = `CIPHERTEXT_WIDTH'd14021333;
cipher_text[8] = `CIPHERTEXT_WIDTH'd11255683;
cipher_text[9] = `CIPHERTEXT_WIDTH'd11323587;
cipher_text[10] = `CIPHERTEXT_WIDTH'd16565208;
cipher_text[11] = `CIPHERTEXT_WIDTH'd14521959;
cipher_text[12] = `CIPHERTEXT_WIDTH'd1064848;
cipher_text[13] = `CIPHERTEXT_WIDTH'd5493216;
cipher_text[14] = `CIPHERTEXT_WIDTH'd12757066;
cipher_text[15] = `CIPHERTEXT_WIDTH'd11483430;
cipher_text[16] = `CIPHERTEXT_WIDTH'd1143571;
cipher_text[17] = `CIPHERTEXT_WIDTH'd3577403;
cipher_text[18] = `CIPHERTEXT_WIDTH'd5348892;
cipher_text[19] = `CIPHERTEXT_WIDTH'd7553633;
cipher_text[20] = `CIPHERTEXT_WIDTH'd2347881;
cipher_text[21] = `CIPHERTEXT_WIDTH'd7512497;
cipher_text[22] = `CIPHERTEXT_WIDTH'd11638147;
cipher_text[23] = `CIPHERTEXT_WIDTH'd11969303;
cipher_text[24] = `CIPHERTEXT_WIDTH'd10308678;
cipher_text[25] = `CIPHERTEXT_WIDTH'd13360669;
cipher_text[26] = `CIPHERTEXT_WIDTH'd10798562;
cipher_text[27] = `CIPHERTEXT_WIDTH'd3677233;
cipher_text[28] = `CIPHERTEXT_WIDTH'd994804;
cipher_text[29] = `CIPHERTEXT_WIDTH'd1059084;
cipher_text[30] = `CIPHERTEXT_WIDTH'd1638275;
cipher_text[31] = `CIPHERTEXT_WIDTH'd8237928;
cipher_text[32] = `CIPHERTEXT_WIDTH'd3892833;
cipher_text[33] = `CIPHERTEXT_WIDTH'd8469088;
cipher_text[34] = `CIPHERTEXT_WIDTH'd12073192;
cipher_text[35] = `CIPHERTEXT_WIDTH'd1119283;
cipher_text[36] = `CIPHERTEXT_WIDTH'd6221787;
cipher_text[37] = `CIPHERTEXT_WIDTH'd13199612;
cipher_text[38] = `CIPHERTEXT_WIDTH'd10958934;
cipher_text[39] = `CIPHERTEXT_WIDTH'd404792;
cipher_text[40] = `CIPHERTEXT_WIDTH'd9420605;
cipher_text[41] = `CIPHERTEXT_WIDTH'd2831257;
cipher_text[42] = `CIPHERTEXT_WIDTH'd11667981;
cipher_text[43] = `CIPHERTEXT_WIDTH'd12437245;
cipher_text[44] = `CIPHERTEXT_WIDTH'd15778611;
cipher_text[45] = `CIPHERTEXT_WIDTH'd6372748;
cipher_text[46] = `CIPHERTEXT_WIDTH'd8499708;
cipher_text[47] = `CIPHERTEXT_WIDTH'd5182833;
cipher_text[48] = `CIPHERTEXT_WIDTH'd15140743;
cipher_text[49] = `CIPHERTEXT_WIDTH'd5332991;
cipher_text[50] = `CIPHERTEXT_WIDTH'd10615171;
cipher_text[51] = `CIPHERTEXT_WIDTH'd9918985;
cipher_text[52] = `CIPHERTEXT_WIDTH'd15739128;
cipher_text[53] = `CIPHERTEXT_WIDTH'd16313453;
cipher_text[54] = `CIPHERTEXT_WIDTH'd10264065;
cipher_text[55] = `CIPHERTEXT_WIDTH'd4107688;
cipher_text[56] = `CIPHERTEXT_WIDTH'd6674337;
cipher_text[57] = `CIPHERTEXT_WIDTH'd6633304;
cipher_text[58] = `CIPHERTEXT_WIDTH'd13717656;
cipher_text[59] = `CIPHERTEXT_WIDTH'd11833555;
cipher_text[60] = `CIPHERTEXT_WIDTH'd7538911;
cipher_text[61] = `CIPHERTEXT_WIDTH'd3814449;
cipher_text[62] = `CIPHERTEXT_WIDTH'd16402355;
cipher_text[63] = `CIPHERTEXT_WIDTH'd3070186;
cipher_text[64] = `CIPHERTEXT_WIDTH'd16636636;
cipher_text[65] = `CIPHERTEXT_WIDTH'd10527559;
cipher_text[66] = `CIPHERTEXT_WIDTH'd13439285;
cipher_text[67] = `CIPHERTEXT_WIDTH'd16225303;
cipher_text[68] = `CIPHERTEXT_WIDTH'd9647030;
cipher_text[69] = `CIPHERTEXT_WIDTH'd1870162;
cipher_text[70] = `CIPHERTEXT_WIDTH'd4328858;
cipher_text[71] = `CIPHERTEXT_WIDTH'd13924049;
cipher_text[72] = `CIPHERTEXT_WIDTH'd5515675;
cipher_text[73] = `CIPHERTEXT_WIDTH'd15239975;
cipher_text[74] = `CIPHERTEXT_WIDTH'd10470506;
cipher_text[75] = `CIPHERTEXT_WIDTH'd2106963;
cipher_text[76] = `CIPHERTEXT_WIDTH'd10783486;
cipher_text[77] = `CIPHERTEXT_WIDTH'd919555;
cipher_text[78] = `CIPHERTEXT_WIDTH'd13520474;
cipher_text[79] = `CIPHERTEXT_WIDTH'd10637024;
cipher_text[80] = `CIPHERTEXT_WIDTH'd3640923;
cipher_text[81] = `CIPHERTEXT_WIDTH'd8149602;
cipher_text[82] = `CIPHERTEXT_WIDTH'd15155742;
cipher_text[83] = `CIPHERTEXT_WIDTH'd2101737;
cipher_text[84] = `CIPHERTEXT_WIDTH'd1814053;
cipher_text[85] = `CIPHERTEXT_WIDTH'd4578513;
cipher_text[86] = `CIPHERTEXT_WIDTH'd10449531;
cipher_text[87] = `CIPHERTEXT_WIDTH'd12135690;
cipher_text[88] = `CIPHERTEXT_WIDTH'd9120479;
cipher_text[89] = `CIPHERTEXT_WIDTH'd16453970;
cipher_text[90] = `CIPHERTEXT_WIDTH'd1522177;
cipher_text[91] = `CIPHERTEXT_WIDTH'd7229675;
cipher_text[92] = `CIPHERTEXT_WIDTH'd5886822;
cipher_text[93] = `CIPHERTEXT_WIDTH'd6900747;
cipher_text[94] = `CIPHERTEXT_WIDTH'd10945115;
cipher_text[95] = `CIPHERTEXT_WIDTH'd14488387;
cipher_text[96] = `CIPHERTEXT_WIDTH'd12721872;
cipher_text[97] = `CIPHERTEXT_WIDTH'd15529862;
cipher_text[98] = `CIPHERTEXT_WIDTH'd3817078;
cipher_text[99] = `CIPHERTEXT_WIDTH'd5460228;
cipher_text[100] = `CIPHERTEXT_WIDTH'd973300;
cipher_text[101] = `CIPHERTEXT_WIDTH'd15183198;
cipher_text[102] = `CIPHERTEXT_WIDTH'd2972823;
cipher_text[103] = `CIPHERTEXT_WIDTH'd10545408;
cipher_text[104] = `CIPHERTEXT_WIDTH'd3277452;
cipher_text[105] = `CIPHERTEXT_WIDTH'd9670290;
cipher_text[106] = `CIPHERTEXT_WIDTH'd9829438;
cipher_text[107] = `CIPHERTEXT_WIDTH'd3617688;
cipher_text[108] = `CIPHERTEXT_WIDTH'd1908915;
cipher_text[109] = `CIPHERTEXT_WIDTH'd2779500;
cipher_text[110] = `CIPHERTEXT_WIDTH'd15149445;
cipher_text[111] = `CIPHERTEXT_WIDTH'd1457914;
cipher_text[112] = `CIPHERTEXT_WIDTH'd14589291;
cipher_text[113] = `CIPHERTEXT_WIDTH'd2499291;
cipher_text[114] = `CIPHERTEXT_WIDTH'd8086120;
cipher_text[115] = `CIPHERTEXT_WIDTH'd15679800;
cipher_text[116] = `CIPHERTEXT_WIDTH'd12752232;
cipher_text[117] = `CIPHERTEXT_WIDTH'd12085796;
cipher_text[118] = `CIPHERTEXT_WIDTH'd5053709;
cipher_text[119] = `CIPHERTEXT_WIDTH'd1603330;
cipher_text[120] = `CIPHERTEXT_WIDTH'd14555380;
cipher_text[121] = `CIPHERTEXT_WIDTH'd15680932;
cipher_text[122] = `CIPHERTEXT_WIDTH'd180513;
cipher_text[123] = `CIPHERTEXT_WIDTH'd2646590;
cipher_text[124] = `CIPHERTEXT_WIDTH'd2031881;
cipher_text[125] = `CIPHERTEXT_WIDTH'd7598057;
cipher_text[126] = `CIPHERTEXT_WIDTH'd14384610;
cipher_text[127] = `CIPHERTEXT_WIDTH'd5725355;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 23;
cipher_text[0] = `CIPHERTEXT_WIDTH'd11627039;
cipher_text[1] = `CIPHERTEXT_WIDTH'd3728060;
cipher_text[2] = `CIPHERTEXT_WIDTH'd4010327;
cipher_text[3] = `CIPHERTEXT_WIDTH'd11258054;
cipher_text[4] = `CIPHERTEXT_WIDTH'd16679980;
cipher_text[5] = `CIPHERTEXT_WIDTH'd11965529;
cipher_text[6] = `CIPHERTEXT_WIDTH'd4485558;
cipher_text[7] = `CIPHERTEXT_WIDTH'd5171541;
cipher_text[8] = `CIPHERTEXT_WIDTH'd6147199;
cipher_text[9] = `CIPHERTEXT_WIDTH'd7731652;
cipher_text[10] = `CIPHERTEXT_WIDTH'd9710772;
cipher_text[11] = `CIPHERTEXT_WIDTH'd1327168;
cipher_text[12] = `CIPHERTEXT_WIDTH'd3582722;
cipher_text[13] = `CIPHERTEXT_WIDTH'd11631572;
cipher_text[14] = `CIPHERTEXT_WIDTH'd6237858;
cipher_text[15] = `CIPHERTEXT_WIDTH'd2571773;
cipher_text[16] = `CIPHERTEXT_WIDTH'd1692881;
cipher_text[17] = `CIPHERTEXT_WIDTH'd88769;
cipher_text[18] = `CIPHERTEXT_WIDTH'd8520589;
cipher_text[19] = `CIPHERTEXT_WIDTH'd3719814;
cipher_text[20] = `CIPHERTEXT_WIDTH'd348903;
cipher_text[21] = `CIPHERTEXT_WIDTH'd16077081;
cipher_text[22] = `CIPHERTEXT_WIDTH'd7199844;
cipher_text[23] = `CIPHERTEXT_WIDTH'd9504942;
cipher_text[24] = `CIPHERTEXT_WIDTH'd564689;
cipher_text[25] = `CIPHERTEXT_WIDTH'd11193643;
cipher_text[26] = `CIPHERTEXT_WIDTH'd16394359;
cipher_text[27] = `CIPHERTEXT_WIDTH'd4356555;
cipher_text[28] = `CIPHERTEXT_WIDTH'd1745029;
cipher_text[29] = `CIPHERTEXT_WIDTH'd15848280;
cipher_text[30] = `CIPHERTEXT_WIDTH'd1754786;
cipher_text[31] = `CIPHERTEXT_WIDTH'd5034145;
cipher_text[32] = `CIPHERTEXT_WIDTH'd10492995;
cipher_text[33] = `CIPHERTEXT_WIDTH'd13074220;
cipher_text[34] = `CIPHERTEXT_WIDTH'd14538054;
cipher_text[35] = `CIPHERTEXT_WIDTH'd1124199;
cipher_text[36] = `CIPHERTEXT_WIDTH'd16429592;
cipher_text[37] = `CIPHERTEXT_WIDTH'd6401938;
cipher_text[38] = `CIPHERTEXT_WIDTH'd10460951;
cipher_text[39] = `CIPHERTEXT_WIDTH'd15983984;
cipher_text[40] = `CIPHERTEXT_WIDTH'd952673;
cipher_text[41] = `CIPHERTEXT_WIDTH'd392876;
cipher_text[42] = `CIPHERTEXT_WIDTH'd8296724;
cipher_text[43] = `CIPHERTEXT_WIDTH'd12274413;
cipher_text[44] = `CIPHERTEXT_WIDTH'd9897797;
cipher_text[45] = `CIPHERTEXT_WIDTH'd8200270;
cipher_text[46] = `CIPHERTEXT_WIDTH'd9081564;
cipher_text[47] = `CIPHERTEXT_WIDTH'd10796267;
cipher_text[48] = `CIPHERTEXT_WIDTH'd3361445;
cipher_text[49] = `CIPHERTEXT_WIDTH'd8747208;
cipher_text[50] = `CIPHERTEXT_WIDTH'd15664126;
cipher_text[51] = `CIPHERTEXT_WIDTH'd14615711;
cipher_text[52] = `CIPHERTEXT_WIDTH'd9389256;
cipher_text[53] = `CIPHERTEXT_WIDTH'd14850898;
cipher_text[54] = `CIPHERTEXT_WIDTH'd1794560;
cipher_text[55] = `CIPHERTEXT_WIDTH'd2910735;
cipher_text[56] = `CIPHERTEXT_WIDTH'd293262;
cipher_text[57] = `CIPHERTEXT_WIDTH'd10301764;
cipher_text[58] = `CIPHERTEXT_WIDTH'd1852774;
cipher_text[59] = `CIPHERTEXT_WIDTH'd6560394;
cipher_text[60] = `CIPHERTEXT_WIDTH'd8871198;
cipher_text[61] = `CIPHERTEXT_WIDTH'd12897897;
cipher_text[62] = `CIPHERTEXT_WIDTH'd3875666;
cipher_text[63] = `CIPHERTEXT_WIDTH'd1723402;
cipher_text[64] = `CIPHERTEXT_WIDTH'd7329944;
cipher_text[65] = `CIPHERTEXT_WIDTH'd1644125;
cipher_text[66] = `CIPHERTEXT_WIDTH'd3958022;
cipher_text[67] = `CIPHERTEXT_WIDTH'd16084678;
cipher_text[68] = `CIPHERTEXT_WIDTH'd8626768;
cipher_text[69] = `CIPHERTEXT_WIDTH'd8945542;
cipher_text[70] = `CIPHERTEXT_WIDTH'd13039833;
cipher_text[71] = `CIPHERTEXT_WIDTH'd11262251;
cipher_text[72] = `CIPHERTEXT_WIDTH'd5579905;
cipher_text[73] = `CIPHERTEXT_WIDTH'd2216713;
cipher_text[74] = `CIPHERTEXT_WIDTH'd16152222;
cipher_text[75] = `CIPHERTEXT_WIDTH'd8204970;
cipher_text[76] = `CIPHERTEXT_WIDTH'd543290;
cipher_text[77] = `CIPHERTEXT_WIDTH'd4632692;
cipher_text[78] = `CIPHERTEXT_WIDTH'd3024694;
cipher_text[79] = `CIPHERTEXT_WIDTH'd11672578;
cipher_text[80] = `CIPHERTEXT_WIDTH'd4431224;
cipher_text[81] = `CIPHERTEXT_WIDTH'd101040;
cipher_text[82] = `CIPHERTEXT_WIDTH'd2443393;
cipher_text[83] = `CIPHERTEXT_WIDTH'd2690947;
cipher_text[84] = `CIPHERTEXT_WIDTH'd5063543;
cipher_text[85] = `CIPHERTEXT_WIDTH'd7747045;
cipher_text[86] = `CIPHERTEXT_WIDTH'd3982381;
cipher_text[87] = `CIPHERTEXT_WIDTH'd15541421;
cipher_text[88] = `CIPHERTEXT_WIDTH'd14379066;
cipher_text[89] = `CIPHERTEXT_WIDTH'd13071852;
cipher_text[90] = `CIPHERTEXT_WIDTH'd13202735;
cipher_text[91] = `CIPHERTEXT_WIDTH'd9819071;
cipher_text[92] = `CIPHERTEXT_WIDTH'd4938597;
cipher_text[93] = `CIPHERTEXT_WIDTH'd8201775;
cipher_text[94] = `CIPHERTEXT_WIDTH'd3292641;
cipher_text[95] = `CIPHERTEXT_WIDTH'd1298682;
cipher_text[96] = `CIPHERTEXT_WIDTH'd5823968;
cipher_text[97] = `CIPHERTEXT_WIDTH'd14414627;
cipher_text[98] = `CIPHERTEXT_WIDTH'd926255;
cipher_text[99] = `CIPHERTEXT_WIDTH'd1946724;
cipher_text[100] = `CIPHERTEXT_WIDTH'd4776659;
cipher_text[101] = `CIPHERTEXT_WIDTH'd16526307;
cipher_text[102] = `CIPHERTEXT_WIDTH'd1587739;
cipher_text[103] = `CIPHERTEXT_WIDTH'd5903718;
cipher_text[104] = `CIPHERTEXT_WIDTH'd7559099;
cipher_text[105] = `CIPHERTEXT_WIDTH'd904076;
cipher_text[106] = `CIPHERTEXT_WIDTH'd5306451;
cipher_text[107] = `CIPHERTEXT_WIDTH'd14817227;
cipher_text[108] = `CIPHERTEXT_WIDTH'd9645742;
cipher_text[109] = `CIPHERTEXT_WIDTH'd2826066;
cipher_text[110] = `CIPHERTEXT_WIDTH'd10883097;
cipher_text[111] = `CIPHERTEXT_WIDTH'd2788285;
cipher_text[112] = `CIPHERTEXT_WIDTH'd9644785;
cipher_text[113] = `CIPHERTEXT_WIDTH'd4892510;
cipher_text[114] = `CIPHERTEXT_WIDTH'd14380889;
cipher_text[115] = `CIPHERTEXT_WIDTH'd11796901;
cipher_text[116] = `CIPHERTEXT_WIDTH'd7971843;
cipher_text[117] = `CIPHERTEXT_WIDTH'd9992330;
cipher_text[118] = `CIPHERTEXT_WIDTH'd15724551;
cipher_text[119] = `CIPHERTEXT_WIDTH'd16658881;
cipher_text[120] = `CIPHERTEXT_WIDTH'd12624869;
cipher_text[121] = `CIPHERTEXT_WIDTH'd4665984;
cipher_text[122] = `CIPHERTEXT_WIDTH'd1471121;
cipher_text[123] = `CIPHERTEXT_WIDTH'd16280783;
cipher_text[124] = `CIPHERTEXT_WIDTH'd922674;
cipher_text[125] = `CIPHERTEXT_WIDTH'd9631922;
cipher_text[126] = `CIPHERTEXT_WIDTH'd3297212;
cipher_text[127] = `CIPHERTEXT_WIDTH'd7231663;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 24;
cipher_text[0] = `CIPHERTEXT_WIDTH'd6454235;
cipher_text[1] = `CIPHERTEXT_WIDTH'd9347816;
cipher_text[2] = `CIPHERTEXT_WIDTH'd13326724;
cipher_text[3] = `CIPHERTEXT_WIDTH'd15151728;
cipher_text[4] = `CIPHERTEXT_WIDTH'd10344787;
cipher_text[5] = `CIPHERTEXT_WIDTH'd16609203;
cipher_text[6] = `CIPHERTEXT_WIDTH'd13640008;
cipher_text[7] = `CIPHERTEXT_WIDTH'd5627996;
cipher_text[8] = `CIPHERTEXT_WIDTH'd5226795;
cipher_text[9] = `CIPHERTEXT_WIDTH'd9427699;
cipher_text[10] = `CIPHERTEXT_WIDTH'd14395475;
cipher_text[11] = `CIPHERTEXT_WIDTH'd16719860;
cipher_text[12] = `CIPHERTEXT_WIDTH'd8857616;
cipher_text[13] = `CIPHERTEXT_WIDTH'd6135054;
cipher_text[14] = `CIPHERTEXT_WIDTH'd16332052;
cipher_text[15] = `CIPHERTEXT_WIDTH'd14360275;
cipher_text[16] = `CIPHERTEXT_WIDTH'd2158034;
cipher_text[17] = `CIPHERTEXT_WIDTH'd11024728;
cipher_text[18] = `CIPHERTEXT_WIDTH'd12320117;
cipher_text[19] = `CIPHERTEXT_WIDTH'd6924973;
cipher_text[20] = `CIPHERTEXT_WIDTH'd10930792;
cipher_text[21] = `CIPHERTEXT_WIDTH'd9533102;
cipher_text[22] = `CIPHERTEXT_WIDTH'd4319881;
cipher_text[23] = `CIPHERTEXT_WIDTH'd10980700;
cipher_text[24] = `CIPHERTEXT_WIDTH'd3709361;
cipher_text[25] = `CIPHERTEXT_WIDTH'd3273773;
cipher_text[26] = `CIPHERTEXT_WIDTH'd1095071;
cipher_text[27] = `CIPHERTEXT_WIDTH'd2610648;
cipher_text[28] = `CIPHERTEXT_WIDTH'd8158091;
cipher_text[29] = `CIPHERTEXT_WIDTH'd2916298;
cipher_text[30] = `CIPHERTEXT_WIDTH'd3164149;
cipher_text[31] = `CIPHERTEXT_WIDTH'd15193823;
cipher_text[32] = `CIPHERTEXT_WIDTH'd16620927;
cipher_text[33] = `CIPHERTEXT_WIDTH'd12822782;
cipher_text[34] = `CIPHERTEXT_WIDTH'd1097896;
cipher_text[35] = `CIPHERTEXT_WIDTH'd5627123;
cipher_text[36] = `CIPHERTEXT_WIDTH'd1112686;
cipher_text[37] = `CIPHERTEXT_WIDTH'd8557434;
cipher_text[38] = `CIPHERTEXT_WIDTH'd5059619;
cipher_text[39] = `CIPHERTEXT_WIDTH'd6455258;
cipher_text[40] = `CIPHERTEXT_WIDTH'd4030963;
cipher_text[41] = `CIPHERTEXT_WIDTH'd13025782;
cipher_text[42] = `CIPHERTEXT_WIDTH'd13096177;
cipher_text[43] = `CIPHERTEXT_WIDTH'd5420025;
cipher_text[44] = `CIPHERTEXT_WIDTH'd11493489;
cipher_text[45] = `CIPHERTEXT_WIDTH'd1883011;
cipher_text[46] = `CIPHERTEXT_WIDTH'd10709747;
cipher_text[47] = `CIPHERTEXT_WIDTH'd2162849;
cipher_text[48] = `CIPHERTEXT_WIDTH'd13735887;
cipher_text[49] = `CIPHERTEXT_WIDTH'd14977136;
cipher_text[50] = `CIPHERTEXT_WIDTH'd15465595;
cipher_text[51] = `CIPHERTEXT_WIDTH'd6546203;
cipher_text[52] = `CIPHERTEXT_WIDTH'd14069800;
cipher_text[53] = `CIPHERTEXT_WIDTH'd416238;
cipher_text[54] = `CIPHERTEXT_WIDTH'd11634955;
cipher_text[55] = `CIPHERTEXT_WIDTH'd2119842;
cipher_text[56] = `CIPHERTEXT_WIDTH'd4603690;
cipher_text[57] = `CIPHERTEXT_WIDTH'd10351288;
cipher_text[58] = `CIPHERTEXT_WIDTH'd140140;
cipher_text[59] = `CIPHERTEXT_WIDTH'd8058232;
cipher_text[60] = `CIPHERTEXT_WIDTH'd16209948;
cipher_text[61] = `CIPHERTEXT_WIDTH'd7923053;
cipher_text[62] = `CIPHERTEXT_WIDTH'd6518434;
cipher_text[63] = `CIPHERTEXT_WIDTH'd1746774;
cipher_text[64] = `CIPHERTEXT_WIDTH'd15782462;
cipher_text[65] = `CIPHERTEXT_WIDTH'd2365750;
cipher_text[66] = `CIPHERTEXT_WIDTH'd12985853;
cipher_text[67] = `CIPHERTEXT_WIDTH'd2915193;
cipher_text[68] = `CIPHERTEXT_WIDTH'd2499565;
cipher_text[69] = `CIPHERTEXT_WIDTH'd137809;
cipher_text[70] = `CIPHERTEXT_WIDTH'd448937;
cipher_text[71] = `CIPHERTEXT_WIDTH'd1600498;
cipher_text[72] = `CIPHERTEXT_WIDTH'd15317766;
cipher_text[73] = `CIPHERTEXT_WIDTH'd4309795;
cipher_text[74] = `CIPHERTEXT_WIDTH'd4937375;
cipher_text[75] = `CIPHERTEXT_WIDTH'd13341630;
cipher_text[76] = `CIPHERTEXT_WIDTH'd16421040;
cipher_text[77] = `CIPHERTEXT_WIDTH'd8864844;
cipher_text[78] = `CIPHERTEXT_WIDTH'd4998085;
cipher_text[79] = `CIPHERTEXT_WIDTH'd8295951;
cipher_text[80] = `CIPHERTEXT_WIDTH'd12213075;
cipher_text[81] = `CIPHERTEXT_WIDTH'd13645085;
cipher_text[82] = `CIPHERTEXT_WIDTH'd14607393;
cipher_text[83] = `CIPHERTEXT_WIDTH'd3077169;
cipher_text[84] = `CIPHERTEXT_WIDTH'd9451829;
cipher_text[85] = `CIPHERTEXT_WIDTH'd11062562;
cipher_text[86] = `CIPHERTEXT_WIDTH'd3063282;
cipher_text[87] = `CIPHERTEXT_WIDTH'd6454682;
cipher_text[88] = `CIPHERTEXT_WIDTH'd12339400;
cipher_text[89] = `CIPHERTEXT_WIDTH'd13376184;
cipher_text[90] = `CIPHERTEXT_WIDTH'd4097003;
cipher_text[91] = `CIPHERTEXT_WIDTH'd805233;
cipher_text[92] = `CIPHERTEXT_WIDTH'd8345518;
cipher_text[93] = `CIPHERTEXT_WIDTH'd8963481;
cipher_text[94] = `CIPHERTEXT_WIDTH'd3894628;
cipher_text[95] = `CIPHERTEXT_WIDTH'd14023401;
cipher_text[96] = `CIPHERTEXT_WIDTH'd2411729;
cipher_text[97] = `CIPHERTEXT_WIDTH'd11044526;
cipher_text[98] = `CIPHERTEXT_WIDTH'd15724051;
cipher_text[99] = `CIPHERTEXT_WIDTH'd3434428;
cipher_text[100] = `CIPHERTEXT_WIDTH'd5019693;
cipher_text[101] = `CIPHERTEXT_WIDTH'd81374;
cipher_text[102] = `CIPHERTEXT_WIDTH'd6855230;
cipher_text[103] = `CIPHERTEXT_WIDTH'd8410703;
cipher_text[104] = `CIPHERTEXT_WIDTH'd608325;
cipher_text[105] = `CIPHERTEXT_WIDTH'd13693833;
cipher_text[106] = `CIPHERTEXT_WIDTH'd14185116;
cipher_text[107] = `CIPHERTEXT_WIDTH'd3241939;
cipher_text[108] = `CIPHERTEXT_WIDTH'd11246365;
cipher_text[109] = `CIPHERTEXT_WIDTH'd4722756;
cipher_text[110] = `CIPHERTEXT_WIDTH'd5040087;
cipher_text[111] = `CIPHERTEXT_WIDTH'd16415445;
cipher_text[112] = `CIPHERTEXT_WIDTH'd9840258;
cipher_text[113] = `CIPHERTEXT_WIDTH'd3769045;
cipher_text[114] = `CIPHERTEXT_WIDTH'd16156969;
cipher_text[115] = `CIPHERTEXT_WIDTH'd5025001;
cipher_text[116] = `CIPHERTEXT_WIDTH'd16491703;
cipher_text[117] = `CIPHERTEXT_WIDTH'd13001961;
cipher_text[118] = `CIPHERTEXT_WIDTH'd4252427;
cipher_text[119] = `CIPHERTEXT_WIDTH'd15317246;
cipher_text[120] = `CIPHERTEXT_WIDTH'd5878733;
cipher_text[121] = `CIPHERTEXT_WIDTH'd15046310;
cipher_text[122] = `CIPHERTEXT_WIDTH'd12776895;
cipher_text[123] = `CIPHERTEXT_WIDTH'd3420166;
cipher_text[124] = `CIPHERTEXT_WIDTH'd10437348;
cipher_text[125] = `CIPHERTEXT_WIDTH'd16013211;
cipher_text[126] = `CIPHERTEXT_WIDTH'd4083884;
cipher_text[127] = `CIPHERTEXT_WIDTH'd14660775;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 25;
cipher_text[0] = `CIPHERTEXT_WIDTH'd8099285;
cipher_text[1] = `CIPHERTEXT_WIDTH'd3382753;
cipher_text[2] = `CIPHERTEXT_WIDTH'd10009198;
cipher_text[3] = `CIPHERTEXT_WIDTH'd5544950;
cipher_text[4] = `CIPHERTEXT_WIDTH'd2401383;
cipher_text[5] = `CIPHERTEXT_WIDTH'd8677778;
cipher_text[6] = `CIPHERTEXT_WIDTH'd12493811;
cipher_text[7] = `CIPHERTEXT_WIDTH'd6151197;
cipher_text[8] = `CIPHERTEXT_WIDTH'd8524149;
cipher_text[9] = `CIPHERTEXT_WIDTH'd15374620;
cipher_text[10] = `CIPHERTEXT_WIDTH'd8897337;
cipher_text[11] = `CIPHERTEXT_WIDTH'd14998217;
cipher_text[12] = `CIPHERTEXT_WIDTH'd3633013;
cipher_text[13] = `CIPHERTEXT_WIDTH'd8193121;
cipher_text[14] = `CIPHERTEXT_WIDTH'd8417052;
cipher_text[15] = `CIPHERTEXT_WIDTH'd10418777;
cipher_text[16] = `CIPHERTEXT_WIDTH'd9605830;
cipher_text[17] = `CIPHERTEXT_WIDTH'd3724400;
cipher_text[18] = `CIPHERTEXT_WIDTH'd8242464;
cipher_text[19] = `CIPHERTEXT_WIDTH'd13251785;
cipher_text[20] = `CIPHERTEXT_WIDTH'd12730891;
cipher_text[21] = `CIPHERTEXT_WIDTH'd8796027;
cipher_text[22] = `CIPHERTEXT_WIDTH'd1766076;
cipher_text[23] = `CIPHERTEXT_WIDTH'd15497377;
cipher_text[24] = `CIPHERTEXT_WIDTH'd12922660;
cipher_text[25] = `CIPHERTEXT_WIDTH'd6077527;
cipher_text[26] = `CIPHERTEXT_WIDTH'd15522245;
cipher_text[27] = `CIPHERTEXT_WIDTH'd11904996;
cipher_text[28] = `CIPHERTEXT_WIDTH'd13429802;
cipher_text[29] = `CIPHERTEXT_WIDTH'd8467398;
cipher_text[30] = `CIPHERTEXT_WIDTH'd9380075;
cipher_text[31] = `CIPHERTEXT_WIDTH'd7131999;
cipher_text[32] = `CIPHERTEXT_WIDTH'd3413213;
cipher_text[33] = `CIPHERTEXT_WIDTH'd13860596;
cipher_text[34] = `CIPHERTEXT_WIDTH'd12731675;
cipher_text[35] = `CIPHERTEXT_WIDTH'd3761221;
cipher_text[36] = `CIPHERTEXT_WIDTH'd8180480;
cipher_text[37] = `CIPHERTEXT_WIDTH'd13231131;
cipher_text[38] = `CIPHERTEXT_WIDTH'd12237283;
cipher_text[39] = `CIPHERTEXT_WIDTH'd12772772;
cipher_text[40] = `CIPHERTEXT_WIDTH'd13499136;
cipher_text[41] = `CIPHERTEXT_WIDTH'd11927477;
cipher_text[42] = `CIPHERTEXT_WIDTH'd8617074;
cipher_text[43] = `CIPHERTEXT_WIDTH'd8740255;
cipher_text[44] = `CIPHERTEXT_WIDTH'd7859312;
cipher_text[45] = `CIPHERTEXT_WIDTH'd15466823;
cipher_text[46] = `CIPHERTEXT_WIDTH'd4329070;
cipher_text[47] = `CIPHERTEXT_WIDTH'd15290572;
cipher_text[48] = `CIPHERTEXT_WIDTH'd6941729;
cipher_text[49] = `CIPHERTEXT_WIDTH'd3969875;
cipher_text[50] = `CIPHERTEXT_WIDTH'd1121612;
cipher_text[51] = `CIPHERTEXT_WIDTH'd9615719;
cipher_text[52] = `CIPHERTEXT_WIDTH'd7904063;
cipher_text[53] = `CIPHERTEXT_WIDTH'd8333617;
cipher_text[54] = `CIPHERTEXT_WIDTH'd5794747;
cipher_text[55] = `CIPHERTEXT_WIDTH'd15942251;
cipher_text[56] = `CIPHERTEXT_WIDTH'd10258859;
cipher_text[57] = `CIPHERTEXT_WIDTH'd1616525;
cipher_text[58] = `CIPHERTEXT_WIDTH'd7330290;
cipher_text[59] = `CIPHERTEXT_WIDTH'd2638547;
cipher_text[60] = `CIPHERTEXT_WIDTH'd8594641;
cipher_text[61] = `CIPHERTEXT_WIDTH'd12899225;
cipher_text[62] = `CIPHERTEXT_WIDTH'd140543;
cipher_text[63] = `CIPHERTEXT_WIDTH'd10051507;
cipher_text[64] = `CIPHERTEXT_WIDTH'd11791051;
cipher_text[65] = `CIPHERTEXT_WIDTH'd1323011;
cipher_text[66] = `CIPHERTEXT_WIDTH'd10863053;
cipher_text[67] = `CIPHERTEXT_WIDTH'd4989494;
cipher_text[68] = `CIPHERTEXT_WIDTH'd2972603;
cipher_text[69] = `CIPHERTEXT_WIDTH'd10559025;
cipher_text[70] = `CIPHERTEXT_WIDTH'd6044744;
cipher_text[71] = `CIPHERTEXT_WIDTH'd9767471;
cipher_text[72] = `CIPHERTEXT_WIDTH'd6742048;
cipher_text[73] = `CIPHERTEXT_WIDTH'd2313868;
cipher_text[74] = `CIPHERTEXT_WIDTH'd10780693;
cipher_text[75] = `CIPHERTEXT_WIDTH'd8715113;
cipher_text[76] = `CIPHERTEXT_WIDTH'd5834696;
cipher_text[77] = `CIPHERTEXT_WIDTH'd14989092;
cipher_text[78] = `CIPHERTEXT_WIDTH'd10372838;
cipher_text[79] = `CIPHERTEXT_WIDTH'd15913546;
cipher_text[80] = `CIPHERTEXT_WIDTH'd13933723;
cipher_text[81] = `CIPHERTEXT_WIDTH'd7848364;
cipher_text[82] = `CIPHERTEXT_WIDTH'd6874905;
cipher_text[83] = `CIPHERTEXT_WIDTH'd2300787;
cipher_text[84] = `CIPHERTEXT_WIDTH'd6459124;
cipher_text[85] = `CIPHERTEXT_WIDTH'd7573665;
cipher_text[86] = `CIPHERTEXT_WIDTH'd7173108;
cipher_text[87] = `CIPHERTEXT_WIDTH'd12789859;
cipher_text[88] = `CIPHERTEXT_WIDTH'd14875165;
cipher_text[89] = `CIPHERTEXT_WIDTH'd15117982;
cipher_text[90] = `CIPHERTEXT_WIDTH'd14246734;
cipher_text[91] = `CIPHERTEXT_WIDTH'd10694590;
cipher_text[92] = `CIPHERTEXT_WIDTH'd10775125;
cipher_text[93] = `CIPHERTEXT_WIDTH'd11332652;
cipher_text[94] = `CIPHERTEXT_WIDTH'd1822529;
cipher_text[95] = `CIPHERTEXT_WIDTH'd2373157;
cipher_text[96] = `CIPHERTEXT_WIDTH'd8474668;
cipher_text[97] = `CIPHERTEXT_WIDTH'd5996763;
cipher_text[98] = `CIPHERTEXT_WIDTH'd6217911;
cipher_text[99] = `CIPHERTEXT_WIDTH'd9531736;
cipher_text[100] = `CIPHERTEXT_WIDTH'd12603468;
cipher_text[101] = `CIPHERTEXT_WIDTH'd14920083;
cipher_text[102] = `CIPHERTEXT_WIDTH'd10274802;
cipher_text[103] = `CIPHERTEXT_WIDTH'd10980193;
cipher_text[104] = `CIPHERTEXT_WIDTH'd9311182;
cipher_text[105] = `CIPHERTEXT_WIDTH'd10151957;
cipher_text[106] = `CIPHERTEXT_WIDTH'd7975531;
cipher_text[107] = `CIPHERTEXT_WIDTH'd12545034;
cipher_text[108] = `CIPHERTEXT_WIDTH'd11720405;
cipher_text[109] = `CIPHERTEXT_WIDTH'd15286804;
cipher_text[110] = `CIPHERTEXT_WIDTH'd2439576;
cipher_text[111] = `CIPHERTEXT_WIDTH'd10494238;
cipher_text[112] = `CIPHERTEXT_WIDTH'd270748;
cipher_text[113] = `CIPHERTEXT_WIDTH'd4158591;
cipher_text[114] = `CIPHERTEXT_WIDTH'd2599477;
cipher_text[115] = `CIPHERTEXT_WIDTH'd15772758;
cipher_text[116] = `CIPHERTEXT_WIDTH'd7009080;
cipher_text[117] = `CIPHERTEXT_WIDTH'd11315176;
cipher_text[118] = `CIPHERTEXT_WIDTH'd11889944;
cipher_text[119] = `CIPHERTEXT_WIDTH'd10464618;
cipher_text[120] = `CIPHERTEXT_WIDTH'd10627270;
cipher_text[121] = `CIPHERTEXT_WIDTH'd3982671;
cipher_text[122] = `CIPHERTEXT_WIDTH'd11790533;
cipher_text[123] = `CIPHERTEXT_WIDTH'd875966;
cipher_text[124] = `CIPHERTEXT_WIDTH'd13023799;
cipher_text[125] = `CIPHERTEXT_WIDTH'd1153955;
cipher_text[126] = `CIPHERTEXT_WIDTH'd6224797;
cipher_text[127] = `CIPHERTEXT_WIDTH'd1423269;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 26;
cipher_text[0] = `CIPHERTEXT_WIDTH'd14443849;
cipher_text[1] = `CIPHERTEXT_WIDTH'd3411792;
cipher_text[2] = `CIPHERTEXT_WIDTH'd15820581;
cipher_text[3] = `CIPHERTEXT_WIDTH'd10922373;
cipher_text[4] = `CIPHERTEXT_WIDTH'd16252737;
cipher_text[5] = `CIPHERTEXT_WIDTH'd6683291;
cipher_text[6] = `CIPHERTEXT_WIDTH'd8175305;
cipher_text[7] = `CIPHERTEXT_WIDTH'd7376342;
cipher_text[8] = `CIPHERTEXT_WIDTH'd14172365;
cipher_text[9] = `CIPHERTEXT_WIDTH'd7763859;
cipher_text[10] = `CIPHERTEXT_WIDTH'd2550992;
cipher_text[11] = `CIPHERTEXT_WIDTH'd8679436;
cipher_text[12] = `CIPHERTEXT_WIDTH'd13787120;
cipher_text[13] = `CIPHERTEXT_WIDTH'd2980311;
cipher_text[14] = `CIPHERTEXT_WIDTH'd1619016;
cipher_text[15] = `CIPHERTEXT_WIDTH'd1682240;
cipher_text[16] = `CIPHERTEXT_WIDTH'd10297541;
cipher_text[17] = `CIPHERTEXT_WIDTH'd4766867;
cipher_text[18] = `CIPHERTEXT_WIDTH'd13243005;
cipher_text[19] = `CIPHERTEXT_WIDTH'd12135249;
cipher_text[20] = `CIPHERTEXT_WIDTH'd1274589;
cipher_text[21] = `CIPHERTEXT_WIDTH'd15311432;
cipher_text[22] = `CIPHERTEXT_WIDTH'd12855334;
cipher_text[23] = `CIPHERTEXT_WIDTH'd7005021;
cipher_text[24] = `CIPHERTEXT_WIDTH'd6850605;
cipher_text[25] = `CIPHERTEXT_WIDTH'd2132601;
cipher_text[26] = `CIPHERTEXT_WIDTH'd9031835;
cipher_text[27] = `CIPHERTEXT_WIDTH'd281209;
cipher_text[28] = `CIPHERTEXT_WIDTH'd11842450;
cipher_text[29] = `CIPHERTEXT_WIDTH'd9302795;
cipher_text[30] = `CIPHERTEXT_WIDTH'd12805540;
cipher_text[31] = `CIPHERTEXT_WIDTH'd4675049;
cipher_text[32] = `CIPHERTEXT_WIDTH'd11203285;
cipher_text[33] = `CIPHERTEXT_WIDTH'd13347463;
cipher_text[34] = `CIPHERTEXT_WIDTH'd3336957;
cipher_text[35] = `CIPHERTEXT_WIDTH'd16404244;
cipher_text[36] = `CIPHERTEXT_WIDTH'd13914585;
cipher_text[37] = `CIPHERTEXT_WIDTH'd12481028;
cipher_text[38] = `CIPHERTEXT_WIDTH'd16449774;
cipher_text[39] = `CIPHERTEXT_WIDTH'd6430406;
cipher_text[40] = `CIPHERTEXT_WIDTH'd9503056;
cipher_text[41] = `CIPHERTEXT_WIDTH'd15951058;
cipher_text[42] = `CIPHERTEXT_WIDTH'd1689803;
cipher_text[43] = `CIPHERTEXT_WIDTH'd10843780;
cipher_text[44] = `CIPHERTEXT_WIDTH'd7172056;
cipher_text[45] = `CIPHERTEXT_WIDTH'd9280645;
cipher_text[46] = `CIPHERTEXT_WIDTH'd14793573;
cipher_text[47] = `CIPHERTEXT_WIDTH'd5861195;
cipher_text[48] = `CIPHERTEXT_WIDTH'd2870539;
cipher_text[49] = `CIPHERTEXT_WIDTH'd16150915;
cipher_text[50] = `CIPHERTEXT_WIDTH'd10609764;
cipher_text[51] = `CIPHERTEXT_WIDTH'd244457;
cipher_text[52] = `CIPHERTEXT_WIDTH'd3237144;
cipher_text[53] = `CIPHERTEXT_WIDTH'd8150952;
cipher_text[54] = `CIPHERTEXT_WIDTH'd3535832;
cipher_text[55] = `CIPHERTEXT_WIDTH'd6406621;
cipher_text[56] = `CIPHERTEXT_WIDTH'd1271018;
cipher_text[57] = `CIPHERTEXT_WIDTH'd10756260;
cipher_text[58] = `CIPHERTEXT_WIDTH'd14953539;
cipher_text[59] = `CIPHERTEXT_WIDTH'd1483565;
cipher_text[60] = `CIPHERTEXT_WIDTH'd3685733;
cipher_text[61] = `CIPHERTEXT_WIDTH'd10084920;
cipher_text[62] = `CIPHERTEXT_WIDTH'd8216523;
cipher_text[63] = `CIPHERTEXT_WIDTH'd11237809;
cipher_text[64] = `CIPHERTEXT_WIDTH'd3839643;
cipher_text[65] = `CIPHERTEXT_WIDTH'd6701135;
cipher_text[66] = `CIPHERTEXT_WIDTH'd1045282;
cipher_text[67] = `CIPHERTEXT_WIDTH'd1178347;
cipher_text[68] = `CIPHERTEXT_WIDTH'd16236822;
cipher_text[69] = `CIPHERTEXT_WIDTH'd10161531;
cipher_text[70] = `CIPHERTEXT_WIDTH'd2374696;
cipher_text[71] = `CIPHERTEXT_WIDTH'd10164612;
cipher_text[72] = `CIPHERTEXT_WIDTH'd3589276;
cipher_text[73] = `CIPHERTEXT_WIDTH'd7945421;
cipher_text[74] = `CIPHERTEXT_WIDTH'd3930466;
cipher_text[75] = `CIPHERTEXT_WIDTH'd5698179;
cipher_text[76] = `CIPHERTEXT_WIDTH'd9137121;
cipher_text[77] = `CIPHERTEXT_WIDTH'd13822973;
cipher_text[78] = `CIPHERTEXT_WIDTH'd11092285;
cipher_text[79] = `CIPHERTEXT_WIDTH'd805890;
cipher_text[80] = `CIPHERTEXT_WIDTH'd2599890;
cipher_text[81] = `CIPHERTEXT_WIDTH'd1693705;
cipher_text[82] = `CIPHERTEXT_WIDTH'd4357469;
cipher_text[83] = `CIPHERTEXT_WIDTH'd15401291;
cipher_text[84] = `CIPHERTEXT_WIDTH'd6235152;
cipher_text[85] = `CIPHERTEXT_WIDTH'd7138905;
cipher_text[86] = `CIPHERTEXT_WIDTH'd10608929;
cipher_text[87] = `CIPHERTEXT_WIDTH'd2282677;
cipher_text[88] = `CIPHERTEXT_WIDTH'd10861192;
cipher_text[89] = `CIPHERTEXT_WIDTH'd6006685;
cipher_text[90] = `CIPHERTEXT_WIDTH'd2097228;
cipher_text[91] = `CIPHERTEXT_WIDTH'd1770453;
cipher_text[92] = `CIPHERTEXT_WIDTH'd3629738;
cipher_text[93] = `CIPHERTEXT_WIDTH'd10550374;
cipher_text[94] = `CIPHERTEXT_WIDTH'd13093943;
cipher_text[95] = `CIPHERTEXT_WIDTH'd14593430;
cipher_text[96] = `CIPHERTEXT_WIDTH'd15914692;
cipher_text[97] = `CIPHERTEXT_WIDTH'd10278538;
cipher_text[98] = `CIPHERTEXT_WIDTH'd15479812;
cipher_text[99] = `CIPHERTEXT_WIDTH'd6968075;
cipher_text[100] = `CIPHERTEXT_WIDTH'd16701150;
cipher_text[101] = `CIPHERTEXT_WIDTH'd13942659;
cipher_text[102] = `CIPHERTEXT_WIDTH'd12481882;
cipher_text[103] = `CIPHERTEXT_WIDTH'd10504584;
cipher_text[104] = `CIPHERTEXT_WIDTH'd6947800;
cipher_text[105] = `CIPHERTEXT_WIDTH'd16092723;
cipher_text[106] = `CIPHERTEXT_WIDTH'd15627305;
cipher_text[107] = `CIPHERTEXT_WIDTH'd7645446;
cipher_text[108] = `CIPHERTEXT_WIDTH'd12346821;
cipher_text[109] = `CIPHERTEXT_WIDTH'd7393003;
cipher_text[110] = `CIPHERTEXT_WIDTH'd15883740;
cipher_text[111] = `CIPHERTEXT_WIDTH'd4446320;
cipher_text[112] = `CIPHERTEXT_WIDTH'd4405684;
cipher_text[113] = `CIPHERTEXT_WIDTH'd14909690;
cipher_text[114] = `CIPHERTEXT_WIDTH'd7461960;
cipher_text[115] = `CIPHERTEXT_WIDTH'd12856065;
cipher_text[116] = `CIPHERTEXT_WIDTH'd14791003;
cipher_text[117] = `CIPHERTEXT_WIDTH'd4967420;
cipher_text[118] = `CIPHERTEXT_WIDTH'd8388173;
cipher_text[119] = `CIPHERTEXT_WIDTH'd13017660;
cipher_text[120] = `CIPHERTEXT_WIDTH'd3825833;
cipher_text[121] = `CIPHERTEXT_WIDTH'd14177644;
cipher_text[122] = `CIPHERTEXT_WIDTH'd9695040;
cipher_text[123] = `CIPHERTEXT_WIDTH'd8347620;
cipher_text[124] = `CIPHERTEXT_WIDTH'd1817718;
cipher_text[125] = `CIPHERTEXT_WIDTH'd12296420;
cipher_text[126] = `CIPHERTEXT_WIDTH'd12600994;
cipher_text[127] = `CIPHERTEXT_WIDTH'd12788713;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 27;
cipher_text[0] = `CIPHERTEXT_WIDTH'd5831600;
cipher_text[1] = `CIPHERTEXT_WIDTH'd12381005;
cipher_text[2] = `CIPHERTEXT_WIDTH'd8180430;
cipher_text[3] = `CIPHERTEXT_WIDTH'd12209314;
cipher_text[4] = `CIPHERTEXT_WIDTH'd11673875;
cipher_text[5] = `CIPHERTEXT_WIDTH'd6450626;
cipher_text[6] = `CIPHERTEXT_WIDTH'd16328147;
cipher_text[7] = `CIPHERTEXT_WIDTH'd1705635;
cipher_text[8] = `CIPHERTEXT_WIDTH'd4386758;
cipher_text[9] = `CIPHERTEXT_WIDTH'd10350708;
cipher_text[10] = `CIPHERTEXT_WIDTH'd207560;
cipher_text[11] = `CIPHERTEXT_WIDTH'd15536053;
cipher_text[12] = `CIPHERTEXT_WIDTH'd299824;
cipher_text[13] = `CIPHERTEXT_WIDTH'd3556184;
cipher_text[14] = `CIPHERTEXT_WIDTH'd510298;
cipher_text[15] = `CIPHERTEXT_WIDTH'd6371264;
cipher_text[16] = `CIPHERTEXT_WIDTH'd3073539;
cipher_text[17] = `CIPHERTEXT_WIDTH'd4862482;
cipher_text[18] = `CIPHERTEXT_WIDTH'd2780517;
cipher_text[19] = `CIPHERTEXT_WIDTH'd13579447;
cipher_text[20] = `CIPHERTEXT_WIDTH'd1260106;
cipher_text[21] = `CIPHERTEXT_WIDTH'd7268635;
cipher_text[22] = `CIPHERTEXT_WIDTH'd9153624;
cipher_text[23] = `CIPHERTEXT_WIDTH'd1419061;
cipher_text[24] = `CIPHERTEXT_WIDTH'd8967043;
cipher_text[25] = `CIPHERTEXT_WIDTH'd2813411;
cipher_text[26] = `CIPHERTEXT_WIDTH'd15252729;
cipher_text[27] = `CIPHERTEXT_WIDTH'd14146202;
cipher_text[28] = `CIPHERTEXT_WIDTH'd9321341;
cipher_text[29] = `CIPHERTEXT_WIDTH'd751289;
cipher_text[30] = `CIPHERTEXT_WIDTH'd5311041;
cipher_text[31] = `CIPHERTEXT_WIDTH'd7834775;
cipher_text[32] = `CIPHERTEXT_WIDTH'd12564735;
cipher_text[33] = `CIPHERTEXT_WIDTH'd4562780;
cipher_text[34] = `CIPHERTEXT_WIDTH'd4272802;
cipher_text[35] = `CIPHERTEXT_WIDTH'd2584811;
cipher_text[36] = `CIPHERTEXT_WIDTH'd8876582;
cipher_text[37] = `CIPHERTEXT_WIDTH'd2673513;
cipher_text[38] = `CIPHERTEXT_WIDTH'd3304333;
cipher_text[39] = `CIPHERTEXT_WIDTH'd13567442;
cipher_text[40] = `CIPHERTEXT_WIDTH'd13039821;
cipher_text[41] = `CIPHERTEXT_WIDTH'd15763853;
cipher_text[42] = `CIPHERTEXT_WIDTH'd1046648;
cipher_text[43] = `CIPHERTEXT_WIDTH'd9965965;
cipher_text[44] = `CIPHERTEXT_WIDTH'd7971915;
cipher_text[45] = `CIPHERTEXT_WIDTH'd12052742;
cipher_text[46] = `CIPHERTEXT_WIDTH'd15950163;
cipher_text[47] = `CIPHERTEXT_WIDTH'd5880997;
cipher_text[48] = `CIPHERTEXT_WIDTH'd11732598;
cipher_text[49] = `CIPHERTEXT_WIDTH'd5442805;
cipher_text[50] = `CIPHERTEXT_WIDTH'd3188221;
cipher_text[51] = `CIPHERTEXT_WIDTH'd4930148;
cipher_text[52] = `CIPHERTEXT_WIDTH'd209022;
cipher_text[53] = `CIPHERTEXT_WIDTH'd5974806;
cipher_text[54] = `CIPHERTEXT_WIDTH'd9748402;
cipher_text[55] = `CIPHERTEXT_WIDTH'd9485219;
cipher_text[56] = `CIPHERTEXT_WIDTH'd10054430;
cipher_text[57] = `CIPHERTEXT_WIDTH'd2223377;
cipher_text[58] = `CIPHERTEXT_WIDTH'd14963770;
cipher_text[59] = `CIPHERTEXT_WIDTH'd4853321;
cipher_text[60] = `CIPHERTEXT_WIDTH'd10519327;
cipher_text[61] = `CIPHERTEXT_WIDTH'd5727692;
cipher_text[62] = `CIPHERTEXT_WIDTH'd13720613;
cipher_text[63] = `CIPHERTEXT_WIDTH'd318919;
cipher_text[64] = `CIPHERTEXT_WIDTH'd2638237;
cipher_text[65] = `CIPHERTEXT_WIDTH'd10510724;
cipher_text[66] = `CIPHERTEXT_WIDTH'd663393;
cipher_text[67] = `CIPHERTEXT_WIDTH'd3674238;
cipher_text[68] = `CIPHERTEXT_WIDTH'd4192819;
cipher_text[69] = `CIPHERTEXT_WIDTH'd14715263;
cipher_text[70] = `CIPHERTEXT_WIDTH'd16435879;
cipher_text[71] = `CIPHERTEXT_WIDTH'd4892687;
cipher_text[72] = `CIPHERTEXT_WIDTH'd6155015;
cipher_text[73] = `CIPHERTEXT_WIDTH'd155157;
cipher_text[74] = `CIPHERTEXT_WIDTH'd2928762;
cipher_text[75] = `CIPHERTEXT_WIDTH'd4877265;
cipher_text[76] = `CIPHERTEXT_WIDTH'd14069639;
cipher_text[77] = `CIPHERTEXT_WIDTH'd9060966;
cipher_text[78] = `CIPHERTEXT_WIDTH'd11656364;
cipher_text[79] = `CIPHERTEXT_WIDTH'd4379635;
cipher_text[80] = `CIPHERTEXT_WIDTH'd16476641;
cipher_text[81] = `CIPHERTEXT_WIDTH'd7792690;
cipher_text[82] = `CIPHERTEXT_WIDTH'd5876147;
cipher_text[83] = `CIPHERTEXT_WIDTH'd10655289;
cipher_text[84] = `CIPHERTEXT_WIDTH'd3114447;
cipher_text[85] = `CIPHERTEXT_WIDTH'd11134625;
cipher_text[86] = `CIPHERTEXT_WIDTH'd12961339;
cipher_text[87] = `CIPHERTEXT_WIDTH'd3465339;
cipher_text[88] = `CIPHERTEXT_WIDTH'd12076550;
cipher_text[89] = `CIPHERTEXT_WIDTH'd6120048;
cipher_text[90] = `CIPHERTEXT_WIDTH'd7756067;
cipher_text[91] = `CIPHERTEXT_WIDTH'd4848559;
cipher_text[92] = `CIPHERTEXT_WIDTH'd12998423;
cipher_text[93] = `CIPHERTEXT_WIDTH'd10186612;
cipher_text[94] = `CIPHERTEXT_WIDTH'd13552458;
cipher_text[95] = `CIPHERTEXT_WIDTH'd7353189;
cipher_text[96] = `CIPHERTEXT_WIDTH'd2565569;
cipher_text[97] = `CIPHERTEXT_WIDTH'd9617145;
cipher_text[98] = `CIPHERTEXT_WIDTH'd2754589;
cipher_text[99] = `CIPHERTEXT_WIDTH'd6490321;
cipher_text[100] = `CIPHERTEXT_WIDTH'd15343570;
cipher_text[101] = `CIPHERTEXT_WIDTH'd13285885;
cipher_text[102] = `CIPHERTEXT_WIDTH'd3240449;
cipher_text[103] = `CIPHERTEXT_WIDTH'd5557630;
cipher_text[104] = `CIPHERTEXT_WIDTH'd14102945;
cipher_text[105] = `CIPHERTEXT_WIDTH'd11875348;
cipher_text[106] = `CIPHERTEXT_WIDTH'd15645432;
cipher_text[107] = `CIPHERTEXT_WIDTH'd15017442;
cipher_text[108] = `CIPHERTEXT_WIDTH'd6274948;
cipher_text[109] = `CIPHERTEXT_WIDTH'd4743144;
cipher_text[110] = `CIPHERTEXT_WIDTH'd14381667;
cipher_text[111] = `CIPHERTEXT_WIDTH'd10699087;
cipher_text[112] = `CIPHERTEXT_WIDTH'd15040210;
cipher_text[113] = `CIPHERTEXT_WIDTH'd11831883;
cipher_text[114] = `CIPHERTEXT_WIDTH'd3361094;
cipher_text[115] = `CIPHERTEXT_WIDTH'd9660717;
cipher_text[116] = `CIPHERTEXT_WIDTH'd3656560;
cipher_text[117] = `CIPHERTEXT_WIDTH'd9245859;
cipher_text[118] = `CIPHERTEXT_WIDTH'd6941198;
cipher_text[119] = `CIPHERTEXT_WIDTH'd2522220;
cipher_text[120] = `CIPHERTEXT_WIDTH'd10655976;
cipher_text[121] = `CIPHERTEXT_WIDTH'd2101325;
cipher_text[122] = `CIPHERTEXT_WIDTH'd5652651;
cipher_text[123] = `CIPHERTEXT_WIDTH'd15002993;
cipher_text[124] = `CIPHERTEXT_WIDTH'd1080454;
cipher_text[125] = `CIPHERTEXT_WIDTH'd12891111;
cipher_text[126] = `CIPHERTEXT_WIDTH'd15305440;
cipher_text[127] = `CIPHERTEXT_WIDTH'd11760722;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 28;
cipher_text[0] = `CIPHERTEXT_WIDTH'd6396680;
cipher_text[1] = `CIPHERTEXT_WIDTH'd10331269;
cipher_text[2] = `CIPHERTEXT_WIDTH'd16762772;
cipher_text[3] = `CIPHERTEXT_WIDTH'd10366141;
cipher_text[4] = `CIPHERTEXT_WIDTH'd8265817;
cipher_text[5] = `CIPHERTEXT_WIDTH'd11952629;
cipher_text[6] = `CIPHERTEXT_WIDTH'd6879378;
cipher_text[7] = `CIPHERTEXT_WIDTH'd14057520;
cipher_text[8] = `CIPHERTEXT_WIDTH'd972402;
cipher_text[9] = `CIPHERTEXT_WIDTH'd6543934;
cipher_text[10] = `CIPHERTEXT_WIDTH'd3013377;
cipher_text[11] = `CIPHERTEXT_WIDTH'd15567730;
cipher_text[12] = `CIPHERTEXT_WIDTH'd11196209;
cipher_text[13] = `CIPHERTEXT_WIDTH'd624513;
cipher_text[14] = `CIPHERTEXT_WIDTH'd16223252;
cipher_text[15] = `CIPHERTEXT_WIDTH'd6090104;
cipher_text[16] = `CIPHERTEXT_WIDTH'd1207884;
cipher_text[17] = `CIPHERTEXT_WIDTH'd13469889;
cipher_text[18] = `CIPHERTEXT_WIDTH'd10650290;
cipher_text[19] = `CIPHERTEXT_WIDTH'd13985758;
cipher_text[20] = `CIPHERTEXT_WIDTH'd6350441;
cipher_text[21] = `CIPHERTEXT_WIDTH'd7933171;
cipher_text[22] = `CIPHERTEXT_WIDTH'd4229756;
cipher_text[23] = `CIPHERTEXT_WIDTH'd11007987;
cipher_text[24] = `CIPHERTEXT_WIDTH'd7044781;
cipher_text[25] = `CIPHERTEXT_WIDTH'd12668133;
cipher_text[26] = `CIPHERTEXT_WIDTH'd16124389;
cipher_text[27] = `CIPHERTEXT_WIDTH'd10833034;
cipher_text[28] = `CIPHERTEXT_WIDTH'd1339249;
cipher_text[29] = `CIPHERTEXT_WIDTH'd3741011;
cipher_text[30] = `CIPHERTEXT_WIDTH'd2963649;
cipher_text[31] = `CIPHERTEXT_WIDTH'd778767;
cipher_text[32] = `CIPHERTEXT_WIDTH'd2876133;
cipher_text[33] = `CIPHERTEXT_WIDTH'd10885734;
cipher_text[34] = `CIPHERTEXT_WIDTH'd10770935;
cipher_text[35] = `CIPHERTEXT_WIDTH'd4976698;
cipher_text[36] = `CIPHERTEXT_WIDTH'd14179131;
cipher_text[37] = `CIPHERTEXT_WIDTH'd4228558;
cipher_text[38] = `CIPHERTEXT_WIDTH'd12595626;
cipher_text[39] = `CIPHERTEXT_WIDTH'd9142103;
cipher_text[40] = `CIPHERTEXT_WIDTH'd9915313;
cipher_text[41] = `CIPHERTEXT_WIDTH'd2692963;
cipher_text[42] = `CIPHERTEXT_WIDTH'd6191159;
cipher_text[43] = `CIPHERTEXT_WIDTH'd261839;
cipher_text[44] = `CIPHERTEXT_WIDTH'd9865208;
cipher_text[45] = `CIPHERTEXT_WIDTH'd10064807;
cipher_text[46] = `CIPHERTEXT_WIDTH'd16444702;
cipher_text[47] = `CIPHERTEXT_WIDTH'd2716271;
cipher_text[48] = `CIPHERTEXT_WIDTH'd5656422;
cipher_text[49] = `CIPHERTEXT_WIDTH'd12061579;
cipher_text[50] = `CIPHERTEXT_WIDTH'd1053486;
cipher_text[51] = `CIPHERTEXT_WIDTH'd13522903;
cipher_text[52] = `CIPHERTEXT_WIDTH'd3910292;
cipher_text[53] = `CIPHERTEXT_WIDTH'd4717340;
cipher_text[54] = `CIPHERTEXT_WIDTH'd11652822;
cipher_text[55] = `CIPHERTEXT_WIDTH'd7551953;
cipher_text[56] = `CIPHERTEXT_WIDTH'd5630492;
cipher_text[57] = `CIPHERTEXT_WIDTH'd11343015;
cipher_text[58] = `CIPHERTEXT_WIDTH'd13132679;
cipher_text[59] = `CIPHERTEXT_WIDTH'd16577948;
cipher_text[60] = `CIPHERTEXT_WIDTH'd16232777;
cipher_text[61] = `CIPHERTEXT_WIDTH'd771619;
cipher_text[62] = `CIPHERTEXT_WIDTH'd16743072;
cipher_text[63] = `CIPHERTEXT_WIDTH'd9589377;
cipher_text[64] = `CIPHERTEXT_WIDTH'd15685913;
cipher_text[65] = `CIPHERTEXT_WIDTH'd996023;
cipher_text[66] = `CIPHERTEXT_WIDTH'd9663711;
cipher_text[67] = `CIPHERTEXT_WIDTH'd2318910;
cipher_text[68] = `CIPHERTEXT_WIDTH'd9172265;
cipher_text[69] = `CIPHERTEXT_WIDTH'd11672889;
cipher_text[70] = `CIPHERTEXT_WIDTH'd14539612;
cipher_text[71] = `CIPHERTEXT_WIDTH'd9987439;
cipher_text[72] = `CIPHERTEXT_WIDTH'd11660413;
cipher_text[73] = `CIPHERTEXT_WIDTH'd4847677;
cipher_text[74] = `CIPHERTEXT_WIDTH'd8073070;
cipher_text[75] = `CIPHERTEXT_WIDTH'd3896609;
cipher_text[76] = `CIPHERTEXT_WIDTH'd2825837;
cipher_text[77] = `CIPHERTEXT_WIDTH'd15375111;
cipher_text[78] = `CIPHERTEXT_WIDTH'd2403248;
cipher_text[79] = `CIPHERTEXT_WIDTH'd12716894;
cipher_text[80] = `CIPHERTEXT_WIDTH'd7046470;
cipher_text[81] = `CIPHERTEXT_WIDTH'd6018470;
cipher_text[82] = `CIPHERTEXT_WIDTH'd11367456;
cipher_text[83] = `CIPHERTEXT_WIDTH'd198252;
cipher_text[84] = `CIPHERTEXT_WIDTH'd11284827;
cipher_text[85] = `CIPHERTEXT_WIDTH'd6817003;
cipher_text[86] = `CIPHERTEXT_WIDTH'd15393549;
cipher_text[87] = `CIPHERTEXT_WIDTH'd16687238;
cipher_text[88] = `CIPHERTEXT_WIDTH'd899412;
cipher_text[89] = `CIPHERTEXT_WIDTH'd7986372;
cipher_text[90] = `CIPHERTEXT_WIDTH'd2497894;
cipher_text[91] = `CIPHERTEXT_WIDTH'd16311272;
cipher_text[92] = `CIPHERTEXT_WIDTH'd381410;
cipher_text[93] = `CIPHERTEXT_WIDTH'd7567057;
cipher_text[94] = `CIPHERTEXT_WIDTH'd7876135;
cipher_text[95] = `CIPHERTEXT_WIDTH'd11797786;
cipher_text[96] = `CIPHERTEXT_WIDTH'd6996715;
cipher_text[97] = `CIPHERTEXT_WIDTH'd8498804;
cipher_text[98] = `CIPHERTEXT_WIDTH'd1353328;
cipher_text[99] = `CIPHERTEXT_WIDTH'd6558038;
cipher_text[100] = `CIPHERTEXT_WIDTH'd10342652;
cipher_text[101] = `CIPHERTEXT_WIDTH'd376070;
cipher_text[102] = `CIPHERTEXT_WIDTH'd3765636;
cipher_text[103] = `CIPHERTEXT_WIDTH'd3621209;
cipher_text[104] = `CIPHERTEXT_WIDTH'd5173757;
cipher_text[105] = `CIPHERTEXT_WIDTH'd10680617;
cipher_text[106] = `CIPHERTEXT_WIDTH'd16328330;
cipher_text[107] = `CIPHERTEXT_WIDTH'd13020737;
cipher_text[108] = `CIPHERTEXT_WIDTH'd16693880;
cipher_text[109] = `CIPHERTEXT_WIDTH'd897895;
cipher_text[110] = `CIPHERTEXT_WIDTH'd3378094;
cipher_text[111] = `CIPHERTEXT_WIDTH'd11995992;
cipher_text[112] = `CIPHERTEXT_WIDTH'd3820033;
cipher_text[113] = `CIPHERTEXT_WIDTH'd1987859;
cipher_text[114] = `CIPHERTEXT_WIDTH'd12575813;
cipher_text[115] = `CIPHERTEXT_WIDTH'd2385375;
cipher_text[116] = `CIPHERTEXT_WIDTH'd603793;
cipher_text[117] = `CIPHERTEXT_WIDTH'd8198888;
cipher_text[118] = `CIPHERTEXT_WIDTH'd5501660;
cipher_text[119] = `CIPHERTEXT_WIDTH'd11853033;
cipher_text[120] = `CIPHERTEXT_WIDTH'd7902237;
cipher_text[121] = `CIPHERTEXT_WIDTH'd4968686;
cipher_text[122] = `CIPHERTEXT_WIDTH'd2290816;
cipher_text[123] = `CIPHERTEXT_WIDTH'd3836739;
cipher_text[124] = `CIPHERTEXT_WIDTH'd7026311;
cipher_text[125] = `CIPHERTEXT_WIDTH'd7151746;
cipher_text[126] = `CIPHERTEXT_WIDTH'd7076429;
cipher_text[127] = `CIPHERTEXT_WIDTH'd15259215;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 29;
cipher_text[0] = `CIPHERTEXT_WIDTH'd16693201;
cipher_text[1] = `CIPHERTEXT_WIDTH'd14192345;
cipher_text[2] = `CIPHERTEXT_WIDTH'd4618013;
cipher_text[3] = `CIPHERTEXT_WIDTH'd13043459;
cipher_text[4] = `CIPHERTEXT_WIDTH'd3766012;
cipher_text[5] = `CIPHERTEXT_WIDTH'd11550177;
cipher_text[6] = `CIPHERTEXT_WIDTH'd6362623;
cipher_text[7] = `CIPHERTEXT_WIDTH'd1628172;
cipher_text[8] = `CIPHERTEXT_WIDTH'd12044122;
cipher_text[9] = `CIPHERTEXT_WIDTH'd3175637;
cipher_text[10] = `CIPHERTEXT_WIDTH'd2064461;
cipher_text[11] = `CIPHERTEXT_WIDTH'd11961323;
cipher_text[12] = `CIPHERTEXT_WIDTH'd8908902;
cipher_text[13] = `CIPHERTEXT_WIDTH'd14927599;
cipher_text[14] = `CIPHERTEXT_WIDTH'd8011961;
cipher_text[15] = `CIPHERTEXT_WIDTH'd9208301;
cipher_text[16] = `CIPHERTEXT_WIDTH'd6368041;
cipher_text[17] = `CIPHERTEXT_WIDTH'd16122038;
cipher_text[18] = `CIPHERTEXT_WIDTH'd8127108;
cipher_text[19] = `CIPHERTEXT_WIDTH'd4702156;
cipher_text[20] = `CIPHERTEXT_WIDTH'd13856271;
cipher_text[21] = `CIPHERTEXT_WIDTH'd9022276;
cipher_text[22] = `CIPHERTEXT_WIDTH'd333098;
cipher_text[23] = `CIPHERTEXT_WIDTH'd977822;
cipher_text[24] = `CIPHERTEXT_WIDTH'd9507370;
cipher_text[25] = `CIPHERTEXT_WIDTH'd8255381;
cipher_text[26] = `CIPHERTEXT_WIDTH'd16410848;
cipher_text[27] = `CIPHERTEXT_WIDTH'd6134652;
cipher_text[28] = `CIPHERTEXT_WIDTH'd4005254;
cipher_text[29] = `CIPHERTEXT_WIDTH'd16095646;
cipher_text[30] = `CIPHERTEXT_WIDTH'd4694164;
cipher_text[31] = `CIPHERTEXT_WIDTH'd720563;
cipher_text[32] = `CIPHERTEXT_WIDTH'd9920517;
cipher_text[33] = `CIPHERTEXT_WIDTH'd14151694;
cipher_text[34] = `CIPHERTEXT_WIDTH'd5239687;
cipher_text[35] = `CIPHERTEXT_WIDTH'd2601137;
cipher_text[36] = `CIPHERTEXT_WIDTH'd10666155;
cipher_text[37] = `CIPHERTEXT_WIDTH'd1164662;
cipher_text[38] = `CIPHERTEXT_WIDTH'd2581555;
cipher_text[39] = `CIPHERTEXT_WIDTH'd7533576;
cipher_text[40] = `CIPHERTEXT_WIDTH'd4391588;
cipher_text[41] = `CIPHERTEXT_WIDTH'd8174069;
cipher_text[42] = `CIPHERTEXT_WIDTH'd13893132;
cipher_text[43] = `CIPHERTEXT_WIDTH'd11887448;
cipher_text[44] = `CIPHERTEXT_WIDTH'd10108760;
cipher_text[45] = `CIPHERTEXT_WIDTH'd14151844;
cipher_text[46] = `CIPHERTEXT_WIDTH'd6007;
cipher_text[47] = `CIPHERTEXT_WIDTH'd3927932;
cipher_text[48] = `CIPHERTEXT_WIDTH'd8148664;
cipher_text[49] = `CIPHERTEXT_WIDTH'd13570499;
cipher_text[50] = `CIPHERTEXT_WIDTH'd6355556;
cipher_text[51] = `CIPHERTEXT_WIDTH'd13014996;
cipher_text[52] = `CIPHERTEXT_WIDTH'd15667618;
cipher_text[53] = `CIPHERTEXT_WIDTH'd3361657;
cipher_text[54] = `CIPHERTEXT_WIDTH'd14056470;
cipher_text[55] = `CIPHERTEXT_WIDTH'd14471922;
cipher_text[56] = `CIPHERTEXT_WIDTH'd1904847;
cipher_text[57] = `CIPHERTEXT_WIDTH'd14471016;
cipher_text[58] = `CIPHERTEXT_WIDTH'd6564674;
cipher_text[59] = `CIPHERTEXT_WIDTH'd12419527;
cipher_text[60] = `CIPHERTEXT_WIDTH'd1258536;
cipher_text[61] = `CIPHERTEXT_WIDTH'd10732708;
cipher_text[62] = `CIPHERTEXT_WIDTH'd1178190;
cipher_text[63] = `CIPHERTEXT_WIDTH'd5199036;
cipher_text[64] = `CIPHERTEXT_WIDTH'd14237608;
cipher_text[65] = `CIPHERTEXT_WIDTH'd3125637;
cipher_text[66] = `CIPHERTEXT_WIDTH'd8321742;
cipher_text[67] = `CIPHERTEXT_WIDTH'd4732696;
cipher_text[68] = `CIPHERTEXT_WIDTH'd1308324;
cipher_text[69] = `CIPHERTEXT_WIDTH'd15016081;
cipher_text[70] = `CIPHERTEXT_WIDTH'd8978096;
cipher_text[71] = `CIPHERTEXT_WIDTH'd10563440;
cipher_text[72] = `CIPHERTEXT_WIDTH'd4460588;
cipher_text[73] = `CIPHERTEXT_WIDTH'd4649605;
cipher_text[74] = `CIPHERTEXT_WIDTH'd14145208;
cipher_text[75] = `CIPHERTEXT_WIDTH'd16463944;
cipher_text[76] = `CIPHERTEXT_WIDTH'd13792953;
cipher_text[77] = `CIPHERTEXT_WIDTH'd9062132;
cipher_text[78] = `CIPHERTEXT_WIDTH'd16162498;
cipher_text[79] = `CIPHERTEXT_WIDTH'd2685651;
cipher_text[80] = `CIPHERTEXT_WIDTH'd1790847;
cipher_text[81] = `CIPHERTEXT_WIDTH'd3471400;
cipher_text[82] = `CIPHERTEXT_WIDTH'd5069701;
cipher_text[83] = `CIPHERTEXT_WIDTH'd9129014;
cipher_text[84] = `CIPHERTEXT_WIDTH'd5221413;
cipher_text[85] = `CIPHERTEXT_WIDTH'd10124191;
cipher_text[86] = `CIPHERTEXT_WIDTH'd6052550;
cipher_text[87] = `CIPHERTEXT_WIDTH'd5129518;
cipher_text[88] = `CIPHERTEXT_WIDTH'd10984496;
cipher_text[89] = `CIPHERTEXT_WIDTH'd13528762;
cipher_text[90] = `CIPHERTEXT_WIDTH'd10281442;
cipher_text[91] = `CIPHERTEXT_WIDTH'd2069731;
cipher_text[92] = `CIPHERTEXT_WIDTH'd14866424;
cipher_text[93] = `CIPHERTEXT_WIDTH'd4967995;
cipher_text[94] = `CIPHERTEXT_WIDTH'd3582605;
cipher_text[95] = `CIPHERTEXT_WIDTH'd7394744;
cipher_text[96] = `CIPHERTEXT_WIDTH'd1785944;
cipher_text[97] = `CIPHERTEXT_WIDTH'd8730088;
cipher_text[98] = `CIPHERTEXT_WIDTH'd14226359;
cipher_text[99] = `CIPHERTEXT_WIDTH'd9933439;
cipher_text[100] = `CIPHERTEXT_WIDTH'd2006355;
cipher_text[101] = `CIPHERTEXT_WIDTH'd8748743;
cipher_text[102] = `CIPHERTEXT_WIDTH'd8130545;
cipher_text[103] = `CIPHERTEXT_WIDTH'd6691507;
cipher_text[104] = `CIPHERTEXT_WIDTH'd11161389;
cipher_text[105] = `CIPHERTEXT_WIDTH'd10704383;
cipher_text[106] = `CIPHERTEXT_WIDTH'd4635552;
cipher_text[107] = `CIPHERTEXT_WIDTH'd2023829;
cipher_text[108] = `CIPHERTEXT_WIDTH'd14090476;
cipher_text[109] = `CIPHERTEXT_WIDTH'd9931146;
cipher_text[110] = `CIPHERTEXT_WIDTH'd15546639;
cipher_text[111] = `CIPHERTEXT_WIDTH'd1859810;
cipher_text[112] = `CIPHERTEXT_WIDTH'd3410232;
cipher_text[113] = `CIPHERTEXT_WIDTH'd16563965;
cipher_text[114] = `CIPHERTEXT_WIDTH'd6271270;
cipher_text[115] = `CIPHERTEXT_WIDTH'd12275632;
cipher_text[116] = `CIPHERTEXT_WIDTH'd3419660;
cipher_text[117] = `CIPHERTEXT_WIDTH'd2202767;
cipher_text[118] = `CIPHERTEXT_WIDTH'd7406756;
cipher_text[119] = `CIPHERTEXT_WIDTH'd14649776;
cipher_text[120] = `CIPHERTEXT_WIDTH'd5096258;
cipher_text[121] = `CIPHERTEXT_WIDTH'd3387550;
cipher_text[122] = `CIPHERTEXT_WIDTH'd3991122;
cipher_text[123] = `CIPHERTEXT_WIDTH'd8871767;
cipher_text[124] = `CIPHERTEXT_WIDTH'd15833297;
cipher_text[125] = `CIPHERTEXT_WIDTH'd4717330;
cipher_text[126] = `CIPHERTEXT_WIDTH'd1159893;
cipher_text[127] = `CIPHERTEXT_WIDTH'd11826224;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 30;
cipher_text[0] = `CIPHERTEXT_WIDTH'd8636805;
cipher_text[1] = `CIPHERTEXT_WIDTH'd8943172;
cipher_text[2] = `CIPHERTEXT_WIDTH'd2635021;
cipher_text[3] = `CIPHERTEXT_WIDTH'd2340977;
cipher_text[4] = `CIPHERTEXT_WIDTH'd15839908;
cipher_text[5] = `CIPHERTEXT_WIDTH'd11371564;
cipher_text[6] = `CIPHERTEXT_WIDTH'd5660276;
cipher_text[7] = `CIPHERTEXT_WIDTH'd633602;
cipher_text[8] = `CIPHERTEXT_WIDTH'd7565422;
cipher_text[9] = `CIPHERTEXT_WIDTH'd13648770;
cipher_text[10] = `CIPHERTEXT_WIDTH'd2097791;
cipher_text[11] = `CIPHERTEXT_WIDTH'd2232167;
cipher_text[12] = `CIPHERTEXT_WIDTH'd1952821;
cipher_text[13] = `CIPHERTEXT_WIDTH'd9262923;
cipher_text[14] = `CIPHERTEXT_WIDTH'd11306843;
cipher_text[15] = `CIPHERTEXT_WIDTH'd31010;
cipher_text[16] = `CIPHERTEXT_WIDTH'd2852236;
cipher_text[17] = `CIPHERTEXT_WIDTH'd6012451;
cipher_text[18] = `CIPHERTEXT_WIDTH'd10449484;
cipher_text[19] = `CIPHERTEXT_WIDTH'd6393495;
cipher_text[20] = `CIPHERTEXT_WIDTH'd2280992;
cipher_text[21] = `CIPHERTEXT_WIDTH'd6230725;
cipher_text[22] = `CIPHERTEXT_WIDTH'd14758385;
cipher_text[23] = `CIPHERTEXT_WIDTH'd3238785;
cipher_text[24] = `CIPHERTEXT_WIDTH'd15414960;
cipher_text[25] = `CIPHERTEXT_WIDTH'd3251497;
cipher_text[26] = `CIPHERTEXT_WIDTH'd11739539;
cipher_text[27] = `CIPHERTEXT_WIDTH'd4530145;
cipher_text[28] = `CIPHERTEXT_WIDTH'd6214853;
cipher_text[29] = `CIPHERTEXT_WIDTH'd2292712;
cipher_text[30] = `CIPHERTEXT_WIDTH'd15153664;
cipher_text[31] = `CIPHERTEXT_WIDTH'd13198147;
cipher_text[32] = `CIPHERTEXT_WIDTH'd9443324;
cipher_text[33] = `CIPHERTEXT_WIDTH'd7988003;
cipher_text[34] = `CIPHERTEXT_WIDTH'd16009377;
cipher_text[35] = `CIPHERTEXT_WIDTH'd7823788;
cipher_text[36] = `CIPHERTEXT_WIDTH'd2123773;
cipher_text[37] = `CIPHERTEXT_WIDTH'd15447479;
cipher_text[38] = `CIPHERTEXT_WIDTH'd2067735;
cipher_text[39] = `CIPHERTEXT_WIDTH'd8468647;
cipher_text[40] = `CIPHERTEXT_WIDTH'd14158996;
cipher_text[41] = `CIPHERTEXT_WIDTH'd2265607;
cipher_text[42] = `CIPHERTEXT_WIDTH'd15140511;
cipher_text[43] = `CIPHERTEXT_WIDTH'd13679766;
cipher_text[44] = `CIPHERTEXT_WIDTH'd11907186;
cipher_text[45] = `CIPHERTEXT_WIDTH'd8998317;
cipher_text[46] = `CIPHERTEXT_WIDTH'd6649826;
cipher_text[47] = `CIPHERTEXT_WIDTH'd15973014;
cipher_text[48] = `CIPHERTEXT_WIDTH'd4227603;
cipher_text[49] = `CIPHERTEXT_WIDTH'd12673642;
cipher_text[50] = `CIPHERTEXT_WIDTH'd8116951;
cipher_text[51] = `CIPHERTEXT_WIDTH'd10363725;
cipher_text[52] = `CIPHERTEXT_WIDTH'd1359282;
cipher_text[53] = `CIPHERTEXT_WIDTH'd13043979;
cipher_text[54] = `CIPHERTEXT_WIDTH'd1738386;
cipher_text[55] = `CIPHERTEXT_WIDTH'd7136476;
cipher_text[56] = `CIPHERTEXT_WIDTH'd13462520;
cipher_text[57] = `CIPHERTEXT_WIDTH'd6314746;
cipher_text[58] = `CIPHERTEXT_WIDTH'd1022607;
cipher_text[59] = `CIPHERTEXT_WIDTH'd7486418;
cipher_text[60] = `CIPHERTEXT_WIDTH'd3302599;
cipher_text[61] = `CIPHERTEXT_WIDTH'd10815847;
cipher_text[62] = `CIPHERTEXT_WIDTH'd2452097;
cipher_text[63] = `CIPHERTEXT_WIDTH'd10578093;
cipher_text[64] = `CIPHERTEXT_WIDTH'd11475960;
cipher_text[65] = `CIPHERTEXT_WIDTH'd5571970;
cipher_text[66] = `CIPHERTEXT_WIDTH'd12217476;
cipher_text[67] = `CIPHERTEXT_WIDTH'd96157;
cipher_text[68] = `CIPHERTEXT_WIDTH'd13129523;
cipher_text[69] = `CIPHERTEXT_WIDTH'd13779049;
cipher_text[70] = `CIPHERTEXT_WIDTH'd4937528;
cipher_text[71] = `CIPHERTEXT_WIDTH'd14406004;
cipher_text[72] = `CIPHERTEXT_WIDTH'd2013886;
cipher_text[73] = `CIPHERTEXT_WIDTH'd9269673;
cipher_text[74] = `CIPHERTEXT_WIDTH'd7701846;
cipher_text[75] = `CIPHERTEXT_WIDTH'd15611827;
cipher_text[76] = `CIPHERTEXT_WIDTH'd11073271;
cipher_text[77] = `CIPHERTEXT_WIDTH'd15447186;
cipher_text[78] = `CIPHERTEXT_WIDTH'd772612;
cipher_text[79] = `CIPHERTEXT_WIDTH'd16320454;
cipher_text[80] = `CIPHERTEXT_WIDTH'd8619059;
cipher_text[81] = `CIPHERTEXT_WIDTH'd13792946;
cipher_text[82] = `CIPHERTEXT_WIDTH'd11740779;
cipher_text[83] = `CIPHERTEXT_WIDTH'd11228740;
cipher_text[84] = `CIPHERTEXT_WIDTH'd6356001;
cipher_text[85] = `CIPHERTEXT_WIDTH'd9963424;
cipher_text[86] = `CIPHERTEXT_WIDTH'd13034656;
cipher_text[87] = `CIPHERTEXT_WIDTH'd12039116;
cipher_text[88] = `CIPHERTEXT_WIDTH'd4166024;
cipher_text[89] = `CIPHERTEXT_WIDTH'd1276902;
cipher_text[90] = `CIPHERTEXT_WIDTH'd6334235;
cipher_text[91] = `CIPHERTEXT_WIDTH'd16149148;
cipher_text[92] = `CIPHERTEXT_WIDTH'd8448863;
cipher_text[93] = `CIPHERTEXT_WIDTH'd5065645;
cipher_text[94] = `CIPHERTEXT_WIDTH'd3267089;
cipher_text[95] = `CIPHERTEXT_WIDTH'd6711272;
cipher_text[96] = `CIPHERTEXT_WIDTH'd5874322;
cipher_text[97] = `CIPHERTEXT_WIDTH'd1937616;
cipher_text[98] = `CIPHERTEXT_WIDTH'd5340914;
cipher_text[99] = `CIPHERTEXT_WIDTH'd16406951;
cipher_text[100] = `CIPHERTEXT_WIDTH'd3905806;
cipher_text[101] = `CIPHERTEXT_WIDTH'd4384425;
cipher_text[102] = `CIPHERTEXT_WIDTH'd13423362;
cipher_text[103] = `CIPHERTEXT_WIDTH'd1983297;
cipher_text[104] = `CIPHERTEXT_WIDTH'd6935813;
cipher_text[105] = `CIPHERTEXT_WIDTH'd8313807;
cipher_text[106] = `CIPHERTEXT_WIDTH'd11496149;
cipher_text[107] = `CIPHERTEXT_WIDTH'd11781058;
cipher_text[108] = `CIPHERTEXT_WIDTH'd6407733;
cipher_text[109] = `CIPHERTEXT_WIDTH'd5745881;
cipher_text[110] = `CIPHERTEXT_WIDTH'd11870267;
cipher_text[111] = `CIPHERTEXT_WIDTH'd199130;
cipher_text[112] = `CIPHERTEXT_WIDTH'd4201511;
cipher_text[113] = `CIPHERTEXT_WIDTH'd1698158;
cipher_text[114] = `CIPHERTEXT_WIDTH'd12433268;
cipher_text[115] = `CIPHERTEXT_WIDTH'd12994965;
cipher_text[116] = `CIPHERTEXT_WIDTH'd5538008;
cipher_text[117] = `CIPHERTEXT_WIDTH'd8884739;
cipher_text[118] = `CIPHERTEXT_WIDTH'd15665314;
cipher_text[119] = `CIPHERTEXT_WIDTH'd5410900;
cipher_text[120] = `CIPHERTEXT_WIDTH'd5783609;
cipher_text[121] = `CIPHERTEXT_WIDTH'd6812272;
cipher_text[122] = `CIPHERTEXT_WIDTH'd8696256;
cipher_text[123] = `CIPHERTEXT_WIDTH'd8960760;
cipher_text[124] = `CIPHERTEXT_WIDTH'd15959764;
cipher_text[125] = `CIPHERTEXT_WIDTH'd5907919;
cipher_text[126] = `CIPHERTEXT_WIDTH'd10118770;
cipher_text[127] = `CIPHERTEXT_WIDTH'd15738757;
rst_n=0;
#100;
rst_n=1;
#100;
row = 0;
skentry = secret_key[0];
ctentry = cipher_text[0];
#20;
row = 1;
skentry = secret_key[1];
ctentry = cipher_text[1];
#20;
row = 2;
skentry = secret_key[2];
ctentry = cipher_text[2];
#20;
row = 3;
skentry = secret_key[3];
ctentry = cipher_text[3];
#20;
row = 4;
skentry = secret_key[4];
ctentry = cipher_text[4];
#20;
row = 5;
skentry = secret_key[5];
ctentry = cipher_text[5];
#20;
row = 6;
skentry = secret_key[6];
ctentry = cipher_text[6];
#20;
row = 7;
skentry = secret_key[7];
ctentry = cipher_text[7];
#20;
row = 8;
skentry = secret_key[8];
ctentry = cipher_text[8];
#20;
row = 9;
skentry = secret_key[9];
ctentry = cipher_text[9];
#20;
row = 10;
skentry = secret_key[10];
ctentry = cipher_text[10];
#20;
row = 11;
skentry = secret_key[11];
ctentry = cipher_text[11];
#20;
row = 12;
skentry = secret_key[12];
ctentry = cipher_text[12];
#20;
row = 13;
skentry = secret_key[13];
ctentry = cipher_text[13];
#20;
row = 14;
skentry = secret_key[14];
ctentry = cipher_text[14];
#20;
row = 15;
skentry = secret_key[15];
ctentry = cipher_text[15];
#20;
row = 16;
skentry = secret_key[16];
ctentry = cipher_text[16];
#20;
row = 17;
skentry = secret_key[17];
ctentry = cipher_text[17];
#20;
row = 18;
skentry = secret_key[18];
ctentry = cipher_text[18];
#20;
row = 19;
skentry = secret_key[19];
ctentry = cipher_text[19];
#20;
row = 20;
skentry = secret_key[20];
ctentry = cipher_text[20];
#20;
row = 21;
skentry = secret_key[21];
ctentry = cipher_text[21];
#20;
row = 22;
skentry = secret_key[22];
ctentry = cipher_text[22];
#20;
row = 23;
skentry = secret_key[23];
ctentry = cipher_text[23];
#20;
row = 24;
skentry = secret_key[24];
ctentry = cipher_text[24];
#20;
row = 25;
skentry = secret_key[25];
ctentry = cipher_text[25];
#20;
row = 26;
skentry = secret_key[26];
ctentry = cipher_text[26];
#20;
row = 27;
skentry = secret_key[27];
ctentry = cipher_text[27];
#20;
row = 28;
skentry = secret_key[28];
ctentry = cipher_text[28];
#20;
row = 29;
skentry = secret_key[29];
ctentry = cipher_text[29];
#20;
row = 30;
skentry = secret_key[30];
ctentry = cipher_text[30];
#20;
row = 31;
skentry = secret_key[31];
ctentry = cipher_text[31];
#20;
row = 32;
skentry = secret_key[32];
ctentry = cipher_text[32];
#20;
row = 33;
skentry = secret_key[33];
ctentry = cipher_text[33];
#20;
row = 34;
skentry = secret_key[34];
ctentry = cipher_text[34];
#20;
row = 35;
skentry = secret_key[35];
ctentry = cipher_text[35];
#20;
row = 36;
skentry = secret_key[36];
ctentry = cipher_text[36];
#20;
row = 37;
skentry = secret_key[37];
ctentry = cipher_text[37];
#20;
row = 38;
skentry = secret_key[38];
ctentry = cipher_text[38];
#20;
row = 39;
skentry = secret_key[39];
ctentry = cipher_text[39];
#20;
row = 40;
skentry = secret_key[40];
ctentry = cipher_text[40];
#20;
row = 41;
skentry = secret_key[41];
ctentry = cipher_text[41];
#20;
row = 42;
skentry = secret_key[42];
ctentry = cipher_text[42];
#20;
row = 43;
skentry = secret_key[43];
ctentry = cipher_text[43];
#20;
row = 44;
skentry = secret_key[44];
ctentry = cipher_text[44];
#20;
row = 45;
skentry = secret_key[45];
ctentry = cipher_text[45];
#20;
row = 46;
skentry = secret_key[46];
ctentry = cipher_text[46];
#20;
row = 47;
skentry = secret_key[47];
ctentry = cipher_text[47];
#20;
row = 48;
skentry = secret_key[48];
ctentry = cipher_text[48];
#20;
row = 49;
skentry = secret_key[49];
ctentry = cipher_text[49];
#20;
row = 50;
skentry = secret_key[50];
ctentry = cipher_text[50];
#20;
row = 51;
skentry = secret_key[51];
ctentry = cipher_text[51];
#20;
row = 52;
skentry = secret_key[52];
ctentry = cipher_text[52];
#20;
row = 53;
skentry = secret_key[53];
ctentry = cipher_text[53];
#20;
row = 54;
skentry = secret_key[54];
ctentry = cipher_text[54];
#20;
row = 55;
skentry = secret_key[55];
ctentry = cipher_text[55];
#20;
row = 56;
skentry = secret_key[56];
ctentry = cipher_text[56];
#20;
row = 57;
skentry = secret_key[57];
ctentry = cipher_text[57];
#20;
row = 58;
skentry = secret_key[58];
ctentry = cipher_text[58];
#20;
row = 59;
skentry = secret_key[59];
ctentry = cipher_text[59];
#20;
row = 60;
skentry = secret_key[60];
ctentry = cipher_text[60];
#20;
row = 61;
skentry = secret_key[61];
ctentry = cipher_text[61];
#20;
row = 62;
skentry = secret_key[62];
ctentry = cipher_text[62];
#20;
row = 63;
skentry = secret_key[63];
ctentry = cipher_text[63];
#20;
row = 64;
skentry = secret_key[64];
ctentry = cipher_text[64];
#20;
row = 65;
skentry = secret_key[65];
ctentry = cipher_text[65];
#20;
row = 66;
skentry = secret_key[66];
ctentry = cipher_text[66];
#20;
row = 67;
skentry = secret_key[67];
ctentry = cipher_text[67];
#20;
row = 68;
skentry = secret_key[68];
ctentry = cipher_text[68];
#20;
row = 69;
skentry = secret_key[69];
ctentry = cipher_text[69];
#20;
row = 70;
skentry = secret_key[70];
ctentry = cipher_text[70];
#20;
row = 71;
skentry = secret_key[71];
ctentry = cipher_text[71];
#20;
row = 72;
skentry = secret_key[72];
ctentry = cipher_text[72];
#20;
row = 73;
skentry = secret_key[73];
ctentry = cipher_text[73];
#20;
row = 74;
skentry = secret_key[74];
ctentry = cipher_text[74];
#20;
row = 75;
skentry = secret_key[75];
ctentry = cipher_text[75];
#20;
row = 76;
skentry = secret_key[76];
ctentry = cipher_text[76];
#20;
row = 77;
skentry = secret_key[77];
ctentry = cipher_text[77];
#20;
row = 78;
skentry = secret_key[78];
ctentry = cipher_text[78];
#20;
row = 79;
skentry = secret_key[79];
ctentry = cipher_text[79];
#20;
row = 80;
skentry = secret_key[80];
ctentry = cipher_text[80];
#20;
row = 81;
skentry = secret_key[81];
ctentry = cipher_text[81];
#20;
row = 82;
skentry = secret_key[82];
ctentry = cipher_text[82];
#20;
row = 83;
skentry = secret_key[83];
ctentry = cipher_text[83];
#20;
row = 84;
skentry = secret_key[84];
ctentry = cipher_text[84];
#20;
row = 85;
skentry = secret_key[85];
ctentry = cipher_text[85];
#20;
row = 86;
skentry = secret_key[86];
ctentry = cipher_text[86];
#20;
row = 87;
skentry = secret_key[87];
ctentry = cipher_text[87];
#20;
row = 88;
skentry = secret_key[88];
ctentry = cipher_text[88];
#20;
row = 89;
skentry = secret_key[89];
ctentry = cipher_text[89];
#20;
row = 90;
skentry = secret_key[90];
ctentry = cipher_text[90];
#20;
row = 91;
skentry = secret_key[91];
ctentry = cipher_text[91];
#20;
row = 92;
skentry = secret_key[92];
ctentry = cipher_text[92];
#20;
row = 93;
skentry = secret_key[93];
ctentry = cipher_text[93];
#20;
row = 94;
skentry = secret_key[94];
ctentry = cipher_text[94];
#20;
row = 95;
skentry = secret_key[95];
ctentry = cipher_text[95];
#20;
row = 96;
skentry = secret_key[96];
ctentry = cipher_text[96];
#20;
row = 97;
skentry = secret_key[97];
ctentry = cipher_text[97];
#20;
row = 98;
skentry = secret_key[98];
ctentry = cipher_text[98];
#20;
row = 99;
skentry = secret_key[99];
ctentry = cipher_text[99];
#20;
row = 100;
skentry = secret_key[100];
ctentry = cipher_text[100];
#20;
row = 101;
skentry = secret_key[101];
ctentry = cipher_text[101];
#20;
row = 102;
skentry = secret_key[102];
ctentry = cipher_text[102];
#20;
row = 103;
skentry = secret_key[103];
ctentry = cipher_text[103];
#20;
row = 104;
skentry = secret_key[104];
ctentry = cipher_text[104];
#20;
row = 105;
skentry = secret_key[105];
ctentry = cipher_text[105];
#20;
row = 106;
skentry = secret_key[106];
ctentry = cipher_text[106];
#20;
row = 107;
skentry = secret_key[107];
ctentry = cipher_text[107];
#20;
row = 108;
skentry = secret_key[108];
ctentry = cipher_text[108];
#20;
row = 109;
skentry = secret_key[109];
ctentry = cipher_text[109];
#20;
row = 110;
skentry = secret_key[110];
ctentry = cipher_text[110];
#20;
row = 111;
skentry = secret_key[111];
ctentry = cipher_text[111];
#20;
row = 112;
skentry = secret_key[112];
ctentry = cipher_text[112];
#20;
row = 113;
skentry = secret_key[113];
ctentry = cipher_text[113];
#20;
row = 114;
skentry = secret_key[114];
ctentry = cipher_text[114];
#20;
row = 115;
skentry = secret_key[115];
ctentry = cipher_text[115];
#20;
row = 116;
skentry = secret_key[116];
ctentry = cipher_text[116];
#20;
row = 117;
skentry = secret_key[117];
ctentry = cipher_text[117];
#20;
row = 118;
skentry = secret_key[118];
ctentry = cipher_text[118];
#20;
row = 119;
skentry = secret_key[119];
ctentry = cipher_text[119];
#20;
row = 120;
skentry = secret_key[120];
ctentry = cipher_text[120];
#20;
row = 121;
skentry = secret_key[121];
ctentry = cipher_text[121];
#20;
row = 122;
skentry = secret_key[122];
ctentry = cipher_text[122];
#20;
row = 123;
skentry = secret_key[123];
ctentry = cipher_text[123];
#20;
row = 124;
skentry = secret_key[124];
ctentry = cipher_text[124];
#20;
row = 125;
skentry = secret_key[125];
ctentry = cipher_text[125];
#20;
row = 126;
skentry = secret_key[126];
ctentry = cipher_text[126];
#20;
row = 127;
skentry = secret_key[127];
ctentry = cipher_text[127];
#20;
$display("Result = %d", result); assert(result == expected);
#20;
expected = 31;
cipher_text[0] = `CIPHERTEXT_WIDTH'd468041;
cipher_text[1] = `CIPHERTEXT_WIDTH'd9101699;
cipher_text[2] = `CIPHERTEXT_WIDTH'd8530744;
cipher_text[3] = `CIPHERTEXT_WIDTH'd12020548;
cipher_text[4] = `CIPHERTEXT_WIDTH'd15952824;
cipher_text[5] = `CIPHERTEXT_WIDTH'd4000422;
cipher_text[6] = `CIPHERTEXT_WIDTH'd7247635;
cipher_text[7] = `CIPHERTEXT_WIDTH'd3694771;
cipher_text[8] = `CIPHERTEXT_WIDTH'd1098332;
cipher_text[9] = `CIPHERTEXT_WIDTH'd720395;
cipher_text[10] = `CIPHERTEXT_WIDTH'd5173570;
cipher_text[11] = `CIPHERTEXT_WIDTH'd16557687;
cipher_text[12] = `CIPHERTEXT_WIDTH'd11913190;
cipher_text[13] = `CIPHERTEXT_WIDTH'd8671251;
cipher_text[14] = `CIPHERTEXT_WIDTH'd5556548;
cipher_text[15] = `CIPHERTEXT_WIDTH'd843405;
cipher_text[16] = `CIPHERTEXT_WIDTH'd9151397;
cipher_text[17] = `CIPHERTEXT_WIDTH'd15739866;
cipher_text[18] = `CIPHERTEXT_WIDTH'd6752991;
cipher_text[19] = `CIPHERTEXT_WIDTH'd5672707;
cipher_text[20] = `CIPHERTEXT_WIDTH'd8286872;
cipher_text[21] = `CIPHERTEXT_WIDTH'd9370370;
cipher_text[22] = `CIPHERTEXT_WIDTH'd15491348;
cipher_text[23] = `CIPHERTEXT_WIDTH'd11750187;
cipher_text[24] = `CIPHERTEXT_WIDTH'd1745023;
cipher_text[25] = `CIPHERTEXT_WIDTH'd8972505;
cipher_text[26] = `CIPHERTEXT_WIDTH'd13428582;
cipher_text[27] = `CIPHERTEXT_WIDTH'd6090856;
cipher_text[28] = `CIPHERTEXT_WIDTH'd3569984;
cipher_text[29] = `CIPHERTEXT_WIDTH'd2437562;
cipher_text[30] = `CIPHERTEXT_WIDTH'd2439384;
cipher_text[31] = `CIPHERTEXT_WIDTH'd10348827;
cipher_text[32] = `CIPHERTEXT_WIDTH'd14458361;
cipher_text[33] = `CIPHERTEXT_WIDTH'd16659254;
cipher_text[34] = `CIPHERTEXT_WIDTH'd10800897;
cipher_text[35] = `CIPHERTEXT_WIDTH'd10948924;
cipher_text[36] = `CIPHERTEXT_WIDTH'd3987541;
cipher_text[37] = `CIPHERTEXT_WIDTH'd12149895;
cipher_text[38] = `CIPHERTEXT_WIDTH'd10300291;
cipher_text[39] = `CIPHERTEXT_WIDTH'd6156729;
cipher_text[40] = `CIPHERTEXT_WIDTH'd14885028;
cipher_text[41] = `CIPHERTEXT_WIDTH'd8790637;
cipher_text[42] = `CIPHERTEXT_WIDTH'd1972374;
cipher_text[43] = `CIPHERTEXT_WIDTH'd2991985;
cipher_text[44] = `CIPHERTEXT_WIDTH'd184607;
cipher_text[45] = `CIPHERTEXT_WIDTH'd12335061;
cipher_text[46] = `CIPHERTEXT_WIDTH'd3872317;
cipher_text[47] = `CIPHERTEXT_WIDTH'd6708592;
cipher_text[48] = `CIPHERTEXT_WIDTH'd15899334;
cipher_text[49] = `CIPHERTEXT_WIDTH'd14641154;
cipher_text[50] = `CIPHERTEXT_WIDTH'd7640778;
cipher_text[51] = `CIPHERTEXT_WIDTH'd6279871;
cipher_text[52] = `CIPHERTEXT_WIDTH'd2493260;
cipher_text[53] = `CIPHERTEXT_WIDTH'd9159512;
cipher_text[54] = `CIPHERTEXT_WIDTH'd8711284;
cipher_text[55] = `CIPHERTEXT_WIDTH'd10616227;
cipher_text[56] = `CIPHERTEXT_WIDTH'd7802758;
cipher_text[57] = `CIPHERTEXT_WIDTH'd16017444;
cipher_text[58] = `CIPHERTEXT_WIDTH'd2500118;
cipher_text[59] = `CIPHERTEXT_WIDTH'd9206650;
cipher_text[60] = `CIPHERTEXT_WIDTH'd3940348;
cipher_text[61] = `CIPHERTEXT_WIDTH'd16043798;
cipher_text[62] = `CIPHERTEXT_WIDTH'd12524808;
cipher_text[63] = `CIPHERTEXT_WIDTH'd9139571;
cipher_text[64] = `CIPHERTEXT_WIDTH'd6696004;
cipher_text[65] = `CIPHERTEXT_WIDTH'd14903309;
cipher_text[66] = `CIPHERTEXT_WIDTH'd263588;
cipher_text[67] = `CIPHERTEXT_WIDTH'd5592951;
cipher_text[68] = `CIPHERTEXT_WIDTH'd8132189;
cipher_text[69] = `CIPHERTEXT_WIDTH'd3324853;
cipher_text[70] = `CIPHERTEXT_WIDTH'd2326950;
cipher_text[71] = `CIPHERTEXT_WIDTH'd5804934;
cipher_text[72] = `CIPHERTEXT_WIDTH'd10008163;
cipher_text[73] = `CIPHERTEXT_WIDTH'd137665;
cipher_text[74] = `CIPHERTEXT_WIDTH'd12042319;
cipher_text[75] = `CIPHERTEXT_WIDTH'd15200290;
cipher_text[76] = `CIPHERTEXT_WIDTH'd2593217;
cipher_text[77] = `CIPHERTEXT_WIDTH'd3020141;
cipher_text[78] = `CIPHERTEXT_WIDTH'd4394509;
cipher_text[79] = `CIPHERTEXT_WIDTH'd14513921;
cipher_text[80] = `CIPHERTEXT_WIDTH'd8044176;
cipher_text[81] = `CIPHERTEXT_WIDTH'd11237050;
cipher_text[82] = `CIPHERTEXT_WIDTH'd9304331;
cipher_text[83] = `CIPHERTEXT_WIDTH'd13504042;
cipher_text[84] = `CIPHERTEXT_WIDTH'd9168041;
cipher_text[85] = `CIPHERTEXT_WIDTH'd3256325;
cipher_text[86] = `CIPHERTEXT_WIDTH'd11543600;
cipher_text[87] = `CIPHERTEXT_WIDTH'd10527861;
cipher_text[88] = `CIPHERTEXT_WIDTH'd7860798;
cipher_text[89] = `CIPHERTEXT_WIDTH'd4904713;
cipher_text[90] = `CIPHERTEXT_WIDTH'd6837191;
cipher_text[91] = `CIPHERTEXT_WIDTH'd9603206;
cipher_text[92] = `CIPHERTEXT_WIDTH'd11587718;
cipher_text[93] = `CIPHERTEXT_WIDTH'd3036512;
cipher_text[94] = `CIPHERTEXT_WIDTH'd6082155;
cipher_text[95] = `CIPHERTEXT_WIDTH'd5379990;
cipher_text[96] = `CIPHERTEXT_WIDTH'd1451676;
cipher_text[97] = `CIPHERTEXT_WIDTH'd4167127;
cipher_text[98] = `CIPHERTEXT_WIDTH'd11330938;
cipher_text[99] = `CIPHERTEXT_WIDTH'd11153274;
cipher_text[100] = `CIPHERTEXT_WIDTH'd15898392;
cipher_text[101] = `CIPHERTEXT_WIDTH'd11051895;
cipher_text[102] = `CIPHERTEXT_WIDTH'd12228177;
cipher_text[103] = `CIPHERTEXT_WIDTH'd7439849;
cipher_text[104] = `CIPHERTEXT_WIDTH'd16474930;
cipher_text[105] = `CIPHERTEXT_WIDTH'd11100493;
cipher_text[106] = `CIPHERTEXT_WIDTH'd16320661;
cipher_text[107] = `CIPHERTEXT_WIDTH'd9363447;
cipher_text[108] = `CIPHERTEXT_WIDTH'd10041706;
cipher_text[109] = `CIPHERTEXT_WIDTH'd1389625;
cipher_text[110] = `CIPHERTEXT_WIDTH'd12457950;
cipher_text[111] = `CIPHERTEXT_WIDTH'd2963777;
cipher_text[112] = `CIPHERTEXT_WIDTH'd16612287;
cipher_text[113] = `CIPHERTEXT_WIDTH'd8756767;
cipher_text[114] = `CIPHERTEXT_WIDTH'd10267416;
cipher_text[115] = `CIPHERTEXT_WIDTH'd5252403;
cipher_text[116] = `CIPHERTEXT_WIDTH'd6876487;
cipher_text[117] = `CIPHERTEXT_WIDTH'd6754220;
cipher_text[118] = `CIPHERTEXT_WIDTH'd3295735;
cipher_text[119] = `CIPHERTEXT_WIDTH'd11388090;
cipher_text[120] = `CIPHERTEXT_WIDTH'd8416602;
cipher_text[121] = `CIPHERTEXT_WIDTH'd12352362;
cipher_text[122] = `CIPHERTEXT_WIDTH'd3981695;
cipher_text[123] = `CIPHERTEXT_WIDTH'd10415450;
cipher_text[124] = `CIPHERTEXT_WIDTH'd8498873;
cipher_text[125] = `CIPHERTEXT_WIDTH'd7201781;
cipher_text[126] = `CIPHERTEXT_WIDTH'd16254597;
cipher_text[127] = `CIPHERTEXT_WIDTH'd6707804;

$finish;
end
endmodule

